module SWCell(
  input  [1:0]  io_q,
  input  [1:0]  io_r,
  input  [15:0] io_e_i,
  input  [15:0] io_f_i,
  input  [15:0] io_ve_i,
  input  [15:0] io_vf_i,
  input  [15:0] io_vv_i,
  output [15:0] io_e_o,
  output [15:0] io_f_o,
  output [15:0] io_v_o
);
  wire [15:0] _T_2 = $signed(io_ve_i) - 16'sh2; // @[SWChisel.scala 78:17]
  wire [15:0] _T_5 = $signed(io_e_i) - 16'sh1; // @[SWChisel.scala 78:39]
  wire [15:0] e_max = $signed(_T_2) >= $signed(_T_5) ? $signed(_T_2) : $signed(_T_5); // @[SWChisel.scala 78:51 79:11 81:11]
  wire [15:0] _T_9 = $signed(io_vf_i) - 16'sh2; // @[SWChisel.scala 85:17]
  wire [15:0] _T_12 = $signed(io_f_i) - 16'sh1; // @[SWChisel.scala 85:38]
  wire [15:0] f_max = $signed(_T_9) > $signed(_T_12) ? $signed(_T_9) : $signed(_T_12); // @[SWChisel.scala 85:50 86:11 88:11]
  wire [15:0] ef_temp = $signed(e_max) > $signed(f_max) ? $signed(e_max) : $signed(f_max); // @[SWChisel.scala 92:24 93:13 95:13]
  wire [15:0] _v_temp_T_2 = $signed(io_vv_i) + 16'sh2; // @[SWChisel.scala 100:23]
  wire [15:0] _v_temp_T_5 = $signed(io_vv_i) - 16'sh2; // @[SWChisel.scala 102:23]
  wire [15:0] v_temp = io_q == io_r ? $signed(_v_temp_T_2) : $signed(_v_temp_T_5); // @[SWChisel.scala 100:12 102:12 99:24]
  assign io_e_o = $signed(_T_2) >= $signed(_T_5) ? $signed(_T_2) : $signed(_T_5); // @[SWChisel.scala 78:51 79:11 81:11]
  assign io_f_o = $signed(_T_9) > $signed(_T_12) ? $signed(_T_9) : $signed(_T_12); // @[SWChisel.scala 85:50 86:11 88:11]
  assign io_v_o = $signed(v_temp) > $signed(ef_temp) ? $signed(v_temp) : $signed(ef_temp); // @[SWChisel.scala 106:27 107:11 109:11]
endmodule
module MyCounter(
  input        clock,
  input        reset,
  input        io_en,
  output [8:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] _io_out_T_2 = io_out + 9'h1; // @[SWChisel.scala 155:55]
  reg [8:0] io_out_r; // @[Reg.scala 35:20]
  assign io_out = io_out_r; // @[SWChisel.scala 155:12]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      io_out_r <= 9'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_out < 9'h190) begin // @[SWChisel.scala 155:28]
        io_out_r <= _io_out_T_2;
      end else begin
        io_out_r <= 9'h0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_out_r = _RAND_0[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MAX(
  input         clock,
  input         reset,
  input         io_start,
  input  [15:0] io_in,
  output        io_done,
  output [15:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] max; // @[SWChisel.scala 122:20]
  reg [8:0] counter; // @[SWChisel.scala 133:24]
  wire [8:0] _counter_T_1 = counter - 9'h1; // @[SWChisel.scala 135:24]
  assign io_done = counter == 9'h0; // @[SWChisel.scala 141:17]
  assign io_out = max; // @[SWChisel.scala 123:10]
  always @(posedge clock) begin
    if (reset) begin // @[SWChisel.scala 122:20]
      max <= 16'sh8000; // @[SWChisel.scala 122:20]
    end else if ($signed(io_in) > $signed(max)) begin // @[SWChisel.scala 126:22]
      max <= io_in; // @[SWChisel.scala 127:9]
    end
    if (reset) begin // @[SWChisel.scala 133:24]
      counter <= 9'h191; // @[SWChisel.scala 133:24]
    end else if (counter == 9'h0) begin // @[SWChisel.scala 141:26]
      counter <= 9'h0; // @[SWChisel.scala 143:13]
    end else if (io_start) begin // @[SWChisel.scala 134:19]
      counter <= _counter_T_1; // @[SWChisel.scala 135:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  max = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SW(
  input         clock,
  input         reset,
  input  [1:0]  io_q_0_b,
  input  [1:0]  io_q_1_b,
  input  [1:0]  io_q_2_b,
  input  [1:0]  io_q_3_b,
  input  [1:0]  io_q_4_b,
  input  [1:0]  io_q_5_b,
  input  [1:0]  io_q_6_b,
  input  [1:0]  io_q_7_b,
  input  [1:0]  io_q_8_b,
  input  [1:0]  io_q_9_b,
  input  [1:0]  io_q_10_b,
  input  [1:0]  io_q_11_b,
  input  [1:0]  io_q_12_b,
  input  [1:0]  io_q_13_b,
  input  [1:0]  io_q_14_b,
  input  [1:0]  io_q_15_b,
  input  [1:0]  io_q_16_b,
  input  [1:0]  io_q_17_b,
  input  [1:0]  io_q_18_b,
  input  [1:0]  io_q_19_b,
  input  [1:0]  io_q_20_b,
  input  [1:0]  io_q_21_b,
  input  [1:0]  io_q_22_b,
  input  [1:0]  io_q_23_b,
  input  [1:0]  io_q_24_b,
  input  [1:0]  io_q_25_b,
  input  [1:0]  io_q_26_b,
  input  [1:0]  io_q_27_b,
  input  [1:0]  io_q_28_b,
  input  [1:0]  io_q_29_b,
  input  [1:0]  io_q_30_b,
  input  [1:0]  io_q_31_b,
  input  [1:0]  io_q_32_b,
  input  [1:0]  io_q_33_b,
  input  [1:0]  io_q_34_b,
  input  [1:0]  io_q_35_b,
  input  [1:0]  io_q_36_b,
  input  [1:0]  io_q_37_b,
  input  [1:0]  io_q_38_b,
  input  [1:0]  io_q_39_b,
  input  [1:0]  io_q_40_b,
  input  [1:0]  io_q_41_b,
  input  [1:0]  io_q_42_b,
  input  [1:0]  io_q_43_b,
  input  [1:0]  io_q_44_b,
  input  [1:0]  io_q_45_b,
  input  [1:0]  io_q_46_b,
  input  [1:0]  io_q_47_b,
  input  [1:0]  io_q_48_b,
  input  [1:0]  io_q_49_b,
  input  [1:0]  io_q_50_b,
  input  [1:0]  io_q_51_b,
  input  [1:0]  io_q_52_b,
  input  [1:0]  io_q_53_b,
  input  [1:0]  io_q_54_b,
  input  [1:0]  io_q_55_b,
  input  [1:0]  io_q_56_b,
  input  [1:0]  io_q_57_b,
  input  [1:0]  io_q_58_b,
  input  [1:0]  io_q_59_b,
  input  [1:0]  io_r_0_b,
  input  [1:0]  io_r_1_b,
  input  [1:0]  io_r_2_b,
  input  [1:0]  io_r_3_b,
  input  [1:0]  io_r_4_b,
  input  [1:0]  io_r_5_b,
  input  [1:0]  io_r_6_b,
  input  [1:0]  io_r_7_b,
  input  [1:0]  io_r_8_b,
  input  [1:0]  io_r_9_b,
  input  [1:0]  io_r_10_b,
  input  [1:0]  io_r_11_b,
  input  [1:0]  io_r_12_b,
  input  [1:0]  io_r_13_b,
  input  [1:0]  io_r_14_b,
  input  [1:0]  io_r_15_b,
  input  [1:0]  io_r_16_b,
  input  [1:0]  io_r_17_b,
  input  [1:0]  io_r_18_b,
  input  [1:0]  io_r_19_b,
  input  [1:0]  io_r_20_b,
  input  [1:0]  io_r_21_b,
  input  [1:0]  io_r_22_b,
  input  [1:0]  io_r_23_b,
  input  [1:0]  io_r_24_b,
  input  [1:0]  io_r_25_b,
  input  [1:0]  io_r_26_b,
  input  [1:0]  io_r_27_b,
  input  [1:0]  io_r_28_b,
  input  [1:0]  io_r_29_b,
  input  [1:0]  io_r_30_b,
  input  [1:0]  io_r_31_b,
  input  [1:0]  io_r_32_b,
  input  [1:0]  io_r_33_b,
  input  [1:0]  io_r_34_b,
  input  [1:0]  io_r_35_b,
  input  [1:0]  io_r_36_b,
  input  [1:0]  io_r_37_b,
  input  [1:0]  io_r_38_b,
  input  [1:0]  io_r_39_b,
  input  [1:0]  io_r_40_b,
  input  [1:0]  io_r_41_b,
  input  [1:0]  io_r_42_b,
  input  [1:0]  io_r_43_b,
  input  [1:0]  io_r_44_b,
  input  [1:0]  io_r_45_b,
  input  [1:0]  io_r_46_b,
  input  [1:0]  io_r_47_b,
  input  [1:0]  io_r_48_b,
  input  [1:0]  io_r_49_b,
  input  [1:0]  io_r_50_b,
  input  [1:0]  io_r_51_b,
  input  [1:0]  io_r_52_b,
  input  [1:0]  io_r_53_b,
  input  [1:0]  io_r_54_b,
  input  [1:0]  io_r_55_b,
  input  [1:0]  io_r_56_b,
  input  [1:0]  io_r_57_b,
  input  [1:0]  io_r_58_b,
  input  [1:0]  io_r_59_b,
  input  [1:0]  io_r_60_b,
  input  [1:0]  io_r_61_b,
  input  [1:0]  io_r_62_b,
  input  [1:0]  io_r_63_b,
  input  [1:0]  io_r_64_b,
  input  [1:0]  io_r_65_b,
  input  [1:0]  io_r_66_b,
  input  [1:0]  io_r_67_b,
  input  [1:0]  io_r_68_b,
  input  [1:0]  io_r_69_b,
  input  [1:0]  io_r_70_b,
  input  [1:0]  io_r_71_b,
  input  [1:0]  io_r_72_b,
  input  [1:0]  io_r_73_b,
  input  [1:0]  io_r_74_b,
  input  [1:0]  io_r_75_b,
  input  [1:0]  io_r_76_b,
  input  [1:0]  io_r_77_b,
  input  [1:0]  io_r_78_b,
  input  [1:0]  io_r_79_b,
  input  [1:0]  io_r_80_b,
  input  [1:0]  io_r_81_b,
  input  [1:0]  io_r_82_b,
  input  [1:0]  io_r_83_b,
  input  [1:0]  io_r_84_b,
  input  [1:0]  io_r_85_b,
  input  [1:0]  io_r_86_b,
  input  [1:0]  io_r_87_b,
  input  [1:0]  io_r_88_b,
  input  [1:0]  io_r_89_b,
  input  [1:0]  io_r_90_b,
  input  [1:0]  io_r_91_b,
  input  [1:0]  io_r_92_b,
  input  [1:0]  io_r_93_b,
  input  [1:0]  io_r_94_b,
  input  [1:0]  io_r_95_b,
  input  [1:0]  io_r_96_b,
  input  [1:0]  io_r_97_b,
  input  [1:0]  io_r_98_b,
  input  [1:0]  io_r_99_b,
  input  [1:0]  io_r_100_b,
  input  [1:0]  io_r_101_b,
  input  [1:0]  io_r_102_b,
  input  [1:0]  io_r_103_b,
  input  [1:0]  io_r_104_b,
  input  [1:0]  io_r_105_b,
  input  [1:0]  io_r_106_b,
  input  [1:0]  io_r_107_b,
  input  [1:0]  io_r_108_b,
  input  [1:0]  io_r_109_b,
  input  [1:0]  io_r_110_b,
  input  [1:0]  io_r_111_b,
  input  [1:0]  io_r_112_b,
  input  [1:0]  io_r_113_b,
  input  [1:0]  io_r_114_b,
  input  [1:0]  io_r_115_b,
  input  [1:0]  io_r_116_b,
  input  [1:0]  io_r_117_b,
  input  [1:0]  io_r_118_b,
  input  [1:0]  io_r_119_b,
  input  [1:0]  io_r_120_b,
  input  [1:0]  io_r_121_b,
  input  [1:0]  io_r_122_b,
  input  [1:0]  io_r_123_b,
  input  [1:0]  io_r_124_b,
  input  [1:0]  io_r_125_b,
  input  [1:0]  io_r_126_b,
  input  [1:0]  io_r_127_b,
  input  [1:0]  io_r_128_b,
  input  [1:0]  io_r_129_b,
  input  [1:0]  io_r_130_b,
  input  [1:0]  io_r_131_b,
  input  [1:0]  io_r_132_b,
  input  [1:0]  io_r_133_b,
  input  [1:0]  io_r_134_b,
  input  [1:0]  io_r_135_b,
  input  [1:0]  io_r_136_b,
  input  [1:0]  io_r_137_b,
  input  [1:0]  io_r_138_b,
  input  [1:0]  io_r_139_b,
  input  [1:0]  io_r_140_b,
  input  [1:0]  io_r_141_b,
  input  [1:0]  io_r_142_b,
  input  [1:0]  io_r_143_b,
  input  [1:0]  io_r_144_b,
  input  [1:0]  io_r_145_b,
  input  [1:0]  io_r_146_b,
  input  [1:0]  io_r_147_b,
  input  [1:0]  io_r_148_b,
  input  [1:0]  io_r_149_b,
  input  [1:0]  io_r_150_b,
  input  [1:0]  io_r_151_b,
  input  [1:0]  io_r_152_b,
  input  [1:0]  io_r_153_b,
  input  [1:0]  io_r_154_b,
  input  [1:0]  io_r_155_b,
  input  [1:0]  io_r_156_b,
  input  [1:0]  io_r_157_b,
  input  [1:0]  io_r_158_b,
  input  [1:0]  io_r_159_b,
  input  [1:0]  io_r_160_b,
  input  [1:0]  io_r_161_b,
  input  [1:0]  io_r_162_b,
  input  [1:0]  io_r_163_b,
  input  [1:0]  io_r_164_b,
  input  [1:0]  io_r_165_b,
  input  [1:0]  io_r_166_b,
  input  [1:0]  io_r_167_b,
  input  [1:0]  io_r_168_b,
  input  [1:0]  io_r_169_b,
  input  [1:0]  io_r_170_b,
  input  [1:0]  io_r_171_b,
  input  [1:0]  io_r_172_b,
  input  [1:0]  io_r_173_b,
  input  [1:0]  io_r_174_b,
  input  [1:0]  io_r_175_b,
  input  [1:0]  io_r_176_b,
  input  [1:0]  io_r_177_b,
  input  [1:0]  io_r_178_b,
  input  [1:0]  io_r_179_b,
  input  [1:0]  io_r_180_b,
  input  [1:0]  io_r_181_b,
  input  [1:0]  io_r_182_b,
  input  [1:0]  io_r_183_b,
  input  [1:0]  io_r_184_b,
  input  [1:0]  io_r_185_b,
  input  [1:0]  io_r_186_b,
  input  [1:0]  io_r_187_b,
  input  [1:0]  io_r_188_b,
  input  [1:0]  io_r_189_b,
  input  [1:0]  io_r_190_b,
  input  [1:0]  io_r_191_b,
  input  [1:0]  io_r_192_b,
  input  [1:0]  io_r_193_b,
  input  [1:0]  io_r_194_b,
  input  [1:0]  io_r_195_b,
  input  [1:0]  io_r_196_b,
  input  [1:0]  io_r_197_b,
  input  [1:0]  io_r_198_b,
  input  [1:0]  io_r_199_b,
  input  [1:0]  io_r_200_b,
  input  [1:0]  io_r_201_b,
  input  [1:0]  io_r_202_b,
  input  [1:0]  io_r_203_b,
  input  [1:0]  io_r_204_b,
  input  [1:0]  io_r_205_b,
  input  [1:0]  io_r_206_b,
  input  [1:0]  io_r_207_b,
  input  [1:0]  io_r_208_b,
  input  [1:0]  io_r_209_b,
  input  [1:0]  io_r_210_b,
  input  [1:0]  io_r_211_b,
  input  [1:0]  io_r_212_b,
  input  [1:0]  io_r_213_b,
  input  [1:0]  io_r_214_b,
  input  [1:0]  io_r_215_b,
  input  [1:0]  io_r_216_b,
  input  [1:0]  io_r_217_b,
  input  [1:0]  io_r_218_b,
  input  [1:0]  io_r_219_b,
  input  [1:0]  io_r_220_b,
  input  [1:0]  io_r_221_b,
  input  [1:0]  io_r_222_b,
  input  [1:0]  io_r_223_b,
  input  [1:0]  io_r_224_b,
  input  [1:0]  io_r_225_b,
  input  [1:0]  io_r_226_b,
  input  [1:0]  io_r_227_b,
  input  [1:0]  io_r_228_b,
  input  [1:0]  io_r_229_b,
  input  [1:0]  io_r_230_b,
  input  [1:0]  io_r_231_b,
  input  [1:0]  io_r_232_b,
  input  [1:0]  io_r_233_b,
  input  [1:0]  io_r_234_b,
  input  [1:0]  io_r_235_b,
  input  [1:0]  io_r_236_b,
  input  [1:0]  io_r_237_b,
  input  [1:0]  io_r_238_b,
  input  [1:0]  io_r_239_b,
  input  [1:0]  io_r_240_b,
  input  [1:0]  io_r_241_b,
  input  [1:0]  io_r_242_b,
  input  [1:0]  io_r_243_b,
  input  [1:0]  io_r_244_b,
  input  [1:0]  io_r_245_b,
  input  [1:0]  io_r_246_b,
  input  [1:0]  io_r_247_b,
  input  [1:0]  io_r_248_b,
  input  [1:0]  io_r_249_b,
  input  [1:0]  io_r_250_b,
  input  [1:0]  io_r_251_b,
  input  [1:0]  io_r_252_b,
  input  [1:0]  io_r_253_b,
  input  [1:0]  io_r_254_b,
  input  [1:0]  io_r_255_b,
  input  [1:0]  io_r_256_b,
  input  [1:0]  io_r_257_b,
  input  [1:0]  io_r_258_b,
  input  [1:0]  io_r_259_b,
  input  [1:0]  io_r_260_b,
  input  [1:0]  io_r_261_b,
  input  [1:0]  io_r_262_b,
  input  [1:0]  io_r_263_b,
  input  [1:0]  io_r_264_b,
  input  [1:0]  io_r_265_b,
  input  [1:0]  io_r_266_b,
  input  [1:0]  io_r_267_b,
  input  [1:0]  io_r_268_b,
  input  [1:0]  io_r_269_b,
  input  [1:0]  io_r_270_b,
  input  [1:0]  io_r_271_b,
  input  [1:0]  io_r_272_b,
  input  [1:0]  io_r_273_b,
  input  [1:0]  io_r_274_b,
  input  [1:0]  io_r_275_b,
  input  [1:0]  io_r_276_b,
  input  [1:0]  io_r_277_b,
  input  [1:0]  io_r_278_b,
  input  [1:0]  io_r_279_b,
  input  [1:0]  io_r_280_b,
  input  [1:0]  io_r_281_b,
  input  [1:0]  io_r_282_b,
  input  [1:0]  io_r_283_b,
  input  [1:0]  io_r_284_b,
  input  [1:0]  io_r_285_b,
  input  [1:0]  io_r_286_b,
  input  [1:0]  io_r_287_b,
  input  [1:0]  io_r_288_b,
  input  [1:0]  io_r_289_b,
  input  [1:0]  io_r_290_b,
  input  [1:0]  io_r_291_b,
  input  [1:0]  io_r_292_b,
  input  [1:0]  io_r_293_b,
  input  [1:0]  io_r_294_b,
  input  [1:0]  io_r_295_b,
  input  [1:0]  io_r_296_b,
  input  [1:0]  io_r_297_b,
  input  [1:0]  io_r_298_b,
  input  [1:0]  io_r_299_b,
  input  [1:0]  io_r_300_b,
  input  [1:0]  io_r_301_b,
  input  [1:0]  io_r_302_b,
  input  [1:0]  io_r_303_b,
  input  [1:0]  io_r_304_b,
  input  [1:0]  io_r_305_b,
  input  [1:0]  io_r_306_b,
  input  [1:0]  io_r_307_b,
  input  [1:0]  io_r_308_b,
  input  [1:0]  io_r_309_b,
  input  [1:0]  io_r_310_b,
  input  [1:0]  io_r_311_b,
  input  [1:0]  io_r_312_b,
  input  [1:0]  io_r_313_b,
  input  [1:0]  io_r_314_b,
  input  [1:0]  io_r_315_b,
  input  [1:0]  io_r_316_b,
  input  [1:0]  io_r_317_b,
  input  [1:0]  io_r_318_b,
  input  [1:0]  io_r_319_b,
  input  [1:0]  io_r_320_b,
  input  [1:0]  io_r_321_b,
  input  [1:0]  io_r_322_b,
  input  [1:0]  io_r_323_b,
  input  [1:0]  io_r_324_b,
  input  [1:0]  io_r_325_b,
  input  [1:0]  io_r_326_b,
  input  [1:0]  io_r_327_b,
  input  [1:0]  io_r_328_b,
  input  [1:0]  io_r_329_b,
  input  [1:0]  io_r_330_b,
  input  [1:0]  io_r_331_b,
  input  [1:0]  io_r_332_b,
  input  [1:0]  io_r_333_b,
  input  [1:0]  io_r_334_b,
  input  [1:0]  io_r_335_b,
  input  [1:0]  io_r_336_b,
  input  [1:0]  io_r_337_b,
  input  [1:0]  io_r_338_b,
  input  [1:0]  io_r_339_b,
  input  [1:0]  io_r_340_b,
  input  [1:0]  io_r_341_b,
  input  [1:0]  io_r_342_b,
  input  [1:0]  io_r_343_b,
  input  [1:0]  io_r_344_b,
  input  [1:0]  io_r_345_b,
  input  [1:0]  io_r_346_b,
  input  [1:0]  io_r_347_b,
  input  [1:0]  io_r_348_b,
  input  [1:0]  io_r_349_b,
  input  [1:0]  io_r_350_b,
  input  [1:0]  io_r_351_b,
  input  [1:0]  io_r_352_b,
  input  [1:0]  io_r_353_b,
  input  [1:0]  io_r_354_b,
  input  [1:0]  io_r_355_b,
  input  [1:0]  io_r_356_b,
  input  [1:0]  io_r_357_b,
  input  [1:0]  io_r_358_b,
  input  [1:0]  io_r_359_b,
  input  [1:0]  io_r_360_b,
  input  [1:0]  io_r_361_b,
  input  [1:0]  io_r_362_b,
  input  [1:0]  io_r_363_b,
  input  [1:0]  io_r_364_b,
  input  [1:0]  io_r_365_b,
  input  [1:0]  io_r_366_b,
  input  [1:0]  io_r_367_b,
  input  [1:0]  io_r_368_b,
  input  [1:0]  io_r_369_b,
  input  [1:0]  io_r_370_b,
  input  [1:0]  io_r_371_b,
  input  [1:0]  io_r_372_b,
  input  [1:0]  io_r_373_b,
  input  [1:0]  io_r_374_b,
  input  [1:0]  io_r_375_b,
  input  [1:0]  io_r_376_b,
  input  [1:0]  io_r_377_b,
  input  [1:0]  io_r_378_b,
  input  [1:0]  io_r_379_b,
  input  [1:0]  io_r_380_b,
  input  [1:0]  io_r_381_b,
  input  [1:0]  io_r_382_b,
  input  [1:0]  io_r_383_b,
  input  [1:0]  io_r_384_b,
  input  [1:0]  io_r_385_b,
  input  [1:0]  io_r_386_b,
  input  [1:0]  io_r_387_b,
  input  [1:0]  io_r_388_b,
  input  [1:0]  io_r_389_b,
  input  [1:0]  io_r_390_b,
  input  [1:0]  io_r_391_b,
  input  [1:0]  io_r_392_b,
  input  [1:0]  io_r_393_b,
  input  [1:0]  io_r_394_b,
  input  [1:0]  io_r_395_b,
  input  [1:0]  io_r_396_b,
  input  [1:0]  io_r_397_b,
  input  [1:0]  io_r_398_b,
  input  [1:0]  io_r_399_b,
  input         io_start,
  output [15:0] io_result,
  output        io_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] array_0_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_0_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_1_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_1_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_2_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_2_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_3_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_3_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_4_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_4_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_5_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_5_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_6_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_6_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_7_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_7_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_8_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_8_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_9_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_9_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_10_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_10_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_11_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_11_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_12_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_12_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_13_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_13_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_14_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_14_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_15_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_15_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_16_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_16_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_17_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_17_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_18_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_18_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_19_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_19_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_20_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_20_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_21_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_21_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_22_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_22_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_23_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_23_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_24_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_24_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_25_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_25_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_26_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_26_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_27_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_27_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_28_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_28_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_29_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_29_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_30_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_30_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_31_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_31_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_32_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_32_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_33_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_33_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_34_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_34_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_35_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_35_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_36_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_36_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_37_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_37_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_38_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_38_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_39_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_39_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_40_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_40_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_41_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_41_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_42_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_42_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_43_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_43_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_44_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_44_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_45_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_45_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_46_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_46_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_47_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_47_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_48_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_48_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_49_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_49_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_50_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_50_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_51_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_51_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_52_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_52_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_53_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_53_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_54_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_54_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_55_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_55_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_56_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_56_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_57_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_57_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_58_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_58_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_59_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_59_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_v_o; // @[SWChisel.scala 170:39]
  wire  r_count_0_clock; // @[SWChisel.scala 171:41]
  wire  r_count_0_reset; // @[SWChisel.scala 171:41]
  wire  r_count_0_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_0_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_1_clock; // @[SWChisel.scala 171:41]
  wire  r_count_1_reset; // @[SWChisel.scala 171:41]
  wire  r_count_1_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_1_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_2_clock; // @[SWChisel.scala 171:41]
  wire  r_count_2_reset; // @[SWChisel.scala 171:41]
  wire  r_count_2_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_2_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_3_clock; // @[SWChisel.scala 171:41]
  wire  r_count_3_reset; // @[SWChisel.scala 171:41]
  wire  r_count_3_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_3_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_4_clock; // @[SWChisel.scala 171:41]
  wire  r_count_4_reset; // @[SWChisel.scala 171:41]
  wire  r_count_4_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_4_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_5_clock; // @[SWChisel.scala 171:41]
  wire  r_count_5_reset; // @[SWChisel.scala 171:41]
  wire  r_count_5_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_5_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_6_clock; // @[SWChisel.scala 171:41]
  wire  r_count_6_reset; // @[SWChisel.scala 171:41]
  wire  r_count_6_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_6_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_7_clock; // @[SWChisel.scala 171:41]
  wire  r_count_7_reset; // @[SWChisel.scala 171:41]
  wire  r_count_7_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_7_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_8_clock; // @[SWChisel.scala 171:41]
  wire  r_count_8_reset; // @[SWChisel.scala 171:41]
  wire  r_count_8_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_8_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_9_clock; // @[SWChisel.scala 171:41]
  wire  r_count_9_reset; // @[SWChisel.scala 171:41]
  wire  r_count_9_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_9_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_10_clock; // @[SWChisel.scala 171:41]
  wire  r_count_10_reset; // @[SWChisel.scala 171:41]
  wire  r_count_10_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_10_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_11_clock; // @[SWChisel.scala 171:41]
  wire  r_count_11_reset; // @[SWChisel.scala 171:41]
  wire  r_count_11_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_11_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_12_clock; // @[SWChisel.scala 171:41]
  wire  r_count_12_reset; // @[SWChisel.scala 171:41]
  wire  r_count_12_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_12_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_13_clock; // @[SWChisel.scala 171:41]
  wire  r_count_13_reset; // @[SWChisel.scala 171:41]
  wire  r_count_13_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_13_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_14_clock; // @[SWChisel.scala 171:41]
  wire  r_count_14_reset; // @[SWChisel.scala 171:41]
  wire  r_count_14_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_14_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_15_clock; // @[SWChisel.scala 171:41]
  wire  r_count_15_reset; // @[SWChisel.scala 171:41]
  wire  r_count_15_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_15_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_16_clock; // @[SWChisel.scala 171:41]
  wire  r_count_16_reset; // @[SWChisel.scala 171:41]
  wire  r_count_16_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_16_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_17_clock; // @[SWChisel.scala 171:41]
  wire  r_count_17_reset; // @[SWChisel.scala 171:41]
  wire  r_count_17_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_17_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_18_clock; // @[SWChisel.scala 171:41]
  wire  r_count_18_reset; // @[SWChisel.scala 171:41]
  wire  r_count_18_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_18_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_19_clock; // @[SWChisel.scala 171:41]
  wire  r_count_19_reset; // @[SWChisel.scala 171:41]
  wire  r_count_19_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_19_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_20_clock; // @[SWChisel.scala 171:41]
  wire  r_count_20_reset; // @[SWChisel.scala 171:41]
  wire  r_count_20_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_20_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_21_clock; // @[SWChisel.scala 171:41]
  wire  r_count_21_reset; // @[SWChisel.scala 171:41]
  wire  r_count_21_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_21_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_22_clock; // @[SWChisel.scala 171:41]
  wire  r_count_22_reset; // @[SWChisel.scala 171:41]
  wire  r_count_22_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_22_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_23_clock; // @[SWChisel.scala 171:41]
  wire  r_count_23_reset; // @[SWChisel.scala 171:41]
  wire  r_count_23_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_23_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_24_clock; // @[SWChisel.scala 171:41]
  wire  r_count_24_reset; // @[SWChisel.scala 171:41]
  wire  r_count_24_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_24_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_25_clock; // @[SWChisel.scala 171:41]
  wire  r_count_25_reset; // @[SWChisel.scala 171:41]
  wire  r_count_25_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_25_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_26_clock; // @[SWChisel.scala 171:41]
  wire  r_count_26_reset; // @[SWChisel.scala 171:41]
  wire  r_count_26_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_26_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_27_clock; // @[SWChisel.scala 171:41]
  wire  r_count_27_reset; // @[SWChisel.scala 171:41]
  wire  r_count_27_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_27_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_28_clock; // @[SWChisel.scala 171:41]
  wire  r_count_28_reset; // @[SWChisel.scala 171:41]
  wire  r_count_28_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_28_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_29_clock; // @[SWChisel.scala 171:41]
  wire  r_count_29_reset; // @[SWChisel.scala 171:41]
  wire  r_count_29_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_29_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_30_clock; // @[SWChisel.scala 171:41]
  wire  r_count_30_reset; // @[SWChisel.scala 171:41]
  wire  r_count_30_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_30_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_31_clock; // @[SWChisel.scala 171:41]
  wire  r_count_31_reset; // @[SWChisel.scala 171:41]
  wire  r_count_31_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_31_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_32_clock; // @[SWChisel.scala 171:41]
  wire  r_count_32_reset; // @[SWChisel.scala 171:41]
  wire  r_count_32_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_32_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_33_clock; // @[SWChisel.scala 171:41]
  wire  r_count_33_reset; // @[SWChisel.scala 171:41]
  wire  r_count_33_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_33_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_34_clock; // @[SWChisel.scala 171:41]
  wire  r_count_34_reset; // @[SWChisel.scala 171:41]
  wire  r_count_34_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_34_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_35_clock; // @[SWChisel.scala 171:41]
  wire  r_count_35_reset; // @[SWChisel.scala 171:41]
  wire  r_count_35_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_35_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_36_clock; // @[SWChisel.scala 171:41]
  wire  r_count_36_reset; // @[SWChisel.scala 171:41]
  wire  r_count_36_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_36_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_37_clock; // @[SWChisel.scala 171:41]
  wire  r_count_37_reset; // @[SWChisel.scala 171:41]
  wire  r_count_37_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_37_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_38_clock; // @[SWChisel.scala 171:41]
  wire  r_count_38_reset; // @[SWChisel.scala 171:41]
  wire  r_count_38_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_38_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_39_clock; // @[SWChisel.scala 171:41]
  wire  r_count_39_reset; // @[SWChisel.scala 171:41]
  wire  r_count_39_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_39_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_40_clock; // @[SWChisel.scala 171:41]
  wire  r_count_40_reset; // @[SWChisel.scala 171:41]
  wire  r_count_40_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_40_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_41_clock; // @[SWChisel.scala 171:41]
  wire  r_count_41_reset; // @[SWChisel.scala 171:41]
  wire  r_count_41_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_41_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_42_clock; // @[SWChisel.scala 171:41]
  wire  r_count_42_reset; // @[SWChisel.scala 171:41]
  wire  r_count_42_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_42_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_43_clock; // @[SWChisel.scala 171:41]
  wire  r_count_43_reset; // @[SWChisel.scala 171:41]
  wire  r_count_43_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_43_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_44_clock; // @[SWChisel.scala 171:41]
  wire  r_count_44_reset; // @[SWChisel.scala 171:41]
  wire  r_count_44_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_44_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_45_clock; // @[SWChisel.scala 171:41]
  wire  r_count_45_reset; // @[SWChisel.scala 171:41]
  wire  r_count_45_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_45_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_46_clock; // @[SWChisel.scala 171:41]
  wire  r_count_46_reset; // @[SWChisel.scala 171:41]
  wire  r_count_46_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_46_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_47_clock; // @[SWChisel.scala 171:41]
  wire  r_count_47_reset; // @[SWChisel.scala 171:41]
  wire  r_count_47_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_47_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_48_clock; // @[SWChisel.scala 171:41]
  wire  r_count_48_reset; // @[SWChisel.scala 171:41]
  wire  r_count_48_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_48_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_49_clock; // @[SWChisel.scala 171:41]
  wire  r_count_49_reset; // @[SWChisel.scala 171:41]
  wire  r_count_49_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_49_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_50_clock; // @[SWChisel.scala 171:41]
  wire  r_count_50_reset; // @[SWChisel.scala 171:41]
  wire  r_count_50_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_50_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_51_clock; // @[SWChisel.scala 171:41]
  wire  r_count_51_reset; // @[SWChisel.scala 171:41]
  wire  r_count_51_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_51_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_52_clock; // @[SWChisel.scala 171:41]
  wire  r_count_52_reset; // @[SWChisel.scala 171:41]
  wire  r_count_52_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_52_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_53_clock; // @[SWChisel.scala 171:41]
  wire  r_count_53_reset; // @[SWChisel.scala 171:41]
  wire  r_count_53_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_53_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_54_clock; // @[SWChisel.scala 171:41]
  wire  r_count_54_reset; // @[SWChisel.scala 171:41]
  wire  r_count_54_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_54_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_55_clock; // @[SWChisel.scala 171:41]
  wire  r_count_55_reset; // @[SWChisel.scala 171:41]
  wire  r_count_55_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_55_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_56_clock; // @[SWChisel.scala 171:41]
  wire  r_count_56_reset; // @[SWChisel.scala 171:41]
  wire  r_count_56_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_56_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_57_clock; // @[SWChisel.scala 171:41]
  wire  r_count_57_reset; // @[SWChisel.scala 171:41]
  wire  r_count_57_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_57_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_58_clock; // @[SWChisel.scala 171:41]
  wire  r_count_58_reset; // @[SWChisel.scala 171:41]
  wire  r_count_58_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_58_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_59_clock; // @[SWChisel.scala 171:41]
  wire  r_count_59_reset; // @[SWChisel.scala 171:41]
  wire  r_count_59_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_59_io_out; // @[SWChisel.scala 171:41]
  wire  max_clock; // @[SWChisel.scala 174:19]
  wire  max_reset; // @[SWChisel.scala 174:19]
  wire  max_io_start; // @[SWChisel.scala 174:19]
  wire [15:0] max_io_in; // @[SWChisel.scala 174:19]
  wire  max_io_done; // @[SWChisel.scala 174:19]
  wire [15:0] max_io_out; // @[SWChisel.scala 174:19]
  reg [15:0] E_0; // @[SWChisel.scala 162:18]
  reg [15:0] E_1; // @[SWChisel.scala 162:18]
  reg [15:0] E_2; // @[SWChisel.scala 162:18]
  reg [15:0] E_3; // @[SWChisel.scala 162:18]
  reg [15:0] E_4; // @[SWChisel.scala 162:18]
  reg [15:0] E_5; // @[SWChisel.scala 162:18]
  reg [15:0] E_6; // @[SWChisel.scala 162:18]
  reg [15:0] E_7; // @[SWChisel.scala 162:18]
  reg [15:0] E_8; // @[SWChisel.scala 162:18]
  reg [15:0] E_9; // @[SWChisel.scala 162:18]
  reg [15:0] E_10; // @[SWChisel.scala 162:18]
  reg [15:0] E_11; // @[SWChisel.scala 162:18]
  reg [15:0] E_12; // @[SWChisel.scala 162:18]
  reg [15:0] E_13; // @[SWChisel.scala 162:18]
  reg [15:0] E_14; // @[SWChisel.scala 162:18]
  reg [15:0] E_15; // @[SWChisel.scala 162:18]
  reg [15:0] E_16; // @[SWChisel.scala 162:18]
  reg [15:0] E_17; // @[SWChisel.scala 162:18]
  reg [15:0] E_18; // @[SWChisel.scala 162:18]
  reg [15:0] E_19; // @[SWChisel.scala 162:18]
  reg [15:0] E_20; // @[SWChisel.scala 162:18]
  reg [15:0] E_21; // @[SWChisel.scala 162:18]
  reg [15:0] E_22; // @[SWChisel.scala 162:18]
  reg [15:0] E_23; // @[SWChisel.scala 162:18]
  reg [15:0] E_24; // @[SWChisel.scala 162:18]
  reg [15:0] E_25; // @[SWChisel.scala 162:18]
  reg [15:0] E_26; // @[SWChisel.scala 162:18]
  reg [15:0] E_27; // @[SWChisel.scala 162:18]
  reg [15:0] E_28; // @[SWChisel.scala 162:18]
  reg [15:0] E_29; // @[SWChisel.scala 162:18]
  reg [15:0] E_30; // @[SWChisel.scala 162:18]
  reg [15:0] E_31; // @[SWChisel.scala 162:18]
  reg [15:0] E_32; // @[SWChisel.scala 162:18]
  reg [15:0] E_33; // @[SWChisel.scala 162:18]
  reg [15:0] E_34; // @[SWChisel.scala 162:18]
  reg [15:0] E_35; // @[SWChisel.scala 162:18]
  reg [15:0] E_36; // @[SWChisel.scala 162:18]
  reg [15:0] E_37; // @[SWChisel.scala 162:18]
  reg [15:0] E_38; // @[SWChisel.scala 162:18]
  reg [15:0] E_39; // @[SWChisel.scala 162:18]
  reg [15:0] E_40; // @[SWChisel.scala 162:18]
  reg [15:0] E_41; // @[SWChisel.scala 162:18]
  reg [15:0] E_42; // @[SWChisel.scala 162:18]
  reg [15:0] E_43; // @[SWChisel.scala 162:18]
  reg [15:0] E_44; // @[SWChisel.scala 162:18]
  reg [15:0] E_45; // @[SWChisel.scala 162:18]
  reg [15:0] E_46; // @[SWChisel.scala 162:18]
  reg [15:0] E_47; // @[SWChisel.scala 162:18]
  reg [15:0] E_48; // @[SWChisel.scala 162:18]
  reg [15:0] E_49; // @[SWChisel.scala 162:18]
  reg [15:0] E_50; // @[SWChisel.scala 162:18]
  reg [15:0] E_51; // @[SWChisel.scala 162:18]
  reg [15:0] E_52; // @[SWChisel.scala 162:18]
  reg [15:0] E_53; // @[SWChisel.scala 162:18]
  reg [15:0] E_54; // @[SWChisel.scala 162:18]
  reg [15:0] E_55; // @[SWChisel.scala 162:18]
  reg [15:0] E_56; // @[SWChisel.scala 162:18]
  reg [15:0] E_57; // @[SWChisel.scala 162:18]
  reg [15:0] E_58; // @[SWChisel.scala 162:18]
  reg [15:0] E_59; // @[SWChisel.scala 162:18]
  reg [15:0] F_1; // @[SWChisel.scala 163:18]
  reg [15:0] F_2; // @[SWChisel.scala 163:18]
  reg [15:0] F_3; // @[SWChisel.scala 163:18]
  reg [15:0] F_4; // @[SWChisel.scala 163:18]
  reg [15:0] F_5; // @[SWChisel.scala 163:18]
  reg [15:0] F_6; // @[SWChisel.scala 163:18]
  reg [15:0] F_7; // @[SWChisel.scala 163:18]
  reg [15:0] F_8; // @[SWChisel.scala 163:18]
  reg [15:0] F_9; // @[SWChisel.scala 163:18]
  reg [15:0] F_10; // @[SWChisel.scala 163:18]
  reg [15:0] F_11; // @[SWChisel.scala 163:18]
  reg [15:0] F_12; // @[SWChisel.scala 163:18]
  reg [15:0] F_13; // @[SWChisel.scala 163:18]
  reg [15:0] F_14; // @[SWChisel.scala 163:18]
  reg [15:0] F_15; // @[SWChisel.scala 163:18]
  reg [15:0] F_16; // @[SWChisel.scala 163:18]
  reg [15:0] F_17; // @[SWChisel.scala 163:18]
  reg [15:0] F_18; // @[SWChisel.scala 163:18]
  reg [15:0] F_19; // @[SWChisel.scala 163:18]
  reg [15:0] F_20; // @[SWChisel.scala 163:18]
  reg [15:0] F_21; // @[SWChisel.scala 163:18]
  reg [15:0] F_22; // @[SWChisel.scala 163:18]
  reg [15:0] F_23; // @[SWChisel.scala 163:18]
  reg [15:0] F_24; // @[SWChisel.scala 163:18]
  reg [15:0] F_25; // @[SWChisel.scala 163:18]
  reg [15:0] F_26; // @[SWChisel.scala 163:18]
  reg [15:0] F_27; // @[SWChisel.scala 163:18]
  reg [15:0] F_28; // @[SWChisel.scala 163:18]
  reg [15:0] F_29; // @[SWChisel.scala 163:18]
  reg [15:0] F_30; // @[SWChisel.scala 163:18]
  reg [15:0] F_31; // @[SWChisel.scala 163:18]
  reg [15:0] F_32; // @[SWChisel.scala 163:18]
  reg [15:0] F_33; // @[SWChisel.scala 163:18]
  reg [15:0] F_34; // @[SWChisel.scala 163:18]
  reg [15:0] F_35; // @[SWChisel.scala 163:18]
  reg [15:0] F_36; // @[SWChisel.scala 163:18]
  reg [15:0] F_37; // @[SWChisel.scala 163:18]
  reg [15:0] F_38; // @[SWChisel.scala 163:18]
  reg [15:0] F_39; // @[SWChisel.scala 163:18]
  reg [15:0] F_40; // @[SWChisel.scala 163:18]
  reg [15:0] F_41; // @[SWChisel.scala 163:18]
  reg [15:0] F_42; // @[SWChisel.scala 163:18]
  reg [15:0] F_43; // @[SWChisel.scala 163:18]
  reg [15:0] F_44; // @[SWChisel.scala 163:18]
  reg [15:0] F_45; // @[SWChisel.scala 163:18]
  reg [15:0] F_46; // @[SWChisel.scala 163:18]
  reg [15:0] F_47; // @[SWChisel.scala 163:18]
  reg [15:0] F_48; // @[SWChisel.scala 163:18]
  reg [15:0] F_49; // @[SWChisel.scala 163:18]
  reg [15:0] F_50; // @[SWChisel.scala 163:18]
  reg [15:0] F_51; // @[SWChisel.scala 163:18]
  reg [15:0] F_52; // @[SWChisel.scala 163:18]
  reg [15:0] F_53; // @[SWChisel.scala 163:18]
  reg [15:0] F_54; // @[SWChisel.scala 163:18]
  reg [15:0] F_55; // @[SWChisel.scala 163:18]
  reg [15:0] F_56; // @[SWChisel.scala 163:18]
  reg [15:0] F_57; // @[SWChisel.scala 163:18]
  reg [15:0] F_58; // @[SWChisel.scala 163:18]
  reg [15:0] F_59; // @[SWChisel.scala 163:18]
  reg [15:0] V1_0; // @[SWChisel.scala 164:19]
  reg [15:0] V1_1; // @[SWChisel.scala 164:19]
  reg [15:0] V1_2; // @[SWChisel.scala 164:19]
  reg [15:0] V1_3; // @[SWChisel.scala 164:19]
  reg [15:0] V1_4; // @[SWChisel.scala 164:19]
  reg [15:0] V1_5; // @[SWChisel.scala 164:19]
  reg [15:0] V1_6; // @[SWChisel.scala 164:19]
  reg [15:0] V1_7; // @[SWChisel.scala 164:19]
  reg [15:0] V1_8; // @[SWChisel.scala 164:19]
  reg [15:0] V1_9; // @[SWChisel.scala 164:19]
  reg [15:0] V1_10; // @[SWChisel.scala 164:19]
  reg [15:0] V1_11; // @[SWChisel.scala 164:19]
  reg [15:0] V1_12; // @[SWChisel.scala 164:19]
  reg [15:0] V1_13; // @[SWChisel.scala 164:19]
  reg [15:0] V1_14; // @[SWChisel.scala 164:19]
  reg [15:0] V1_15; // @[SWChisel.scala 164:19]
  reg [15:0] V1_16; // @[SWChisel.scala 164:19]
  reg [15:0] V1_17; // @[SWChisel.scala 164:19]
  reg [15:0] V1_18; // @[SWChisel.scala 164:19]
  reg [15:0] V1_19; // @[SWChisel.scala 164:19]
  reg [15:0] V1_20; // @[SWChisel.scala 164:19]
  reg [15:0] V1_21; // @[SWChisel.scala 164:19]
  reg [15:0] V1_22; // @[SWChisel.scala 164:19]
  reg [15:0] V1_23; // @[SWChisel.scala 164:19]
  reg [15:0] V1_24; // @[SWChisel.scala 164:19]
  reg [15:0] V1_25; // @[SWChisel.scala 164:19]
  reg [15:0] V1_26; // @[SWChisel.scala 164:19]
  reg [15:0] V1_27; // @[SWChisel.scala 164:19]
  reg [15:0] V1_28; // @[SWChisel.scala 164:19]
  reg [15:0] V1_29; // @[SWChisel.scala 164:19]
  reg [15:0] V1_30; // @[SWChisel.scala 164:19]
  reg [15:0] V1_31; // @[SWChisel.scala 164:19]
  reg [15:0] V1_32; // @[SWChisel.scala 164:19]
  reg [15:0] V1_33; // @[SWChisel.scala 164:19]
  reg [15:0] V1_34; // @[SWChisel.scala 164:19]
  reg [15:0] V1_35; // @[SWChisel.scala 164:19]
  reg [15:0] V1_36; // @[SWChisel.scala 164:19]
  reg [15:0] V1_37; // @[SWChisel.scala 164:19]
  reg [15:0] V1_38; // @[SWChisel.scala 164:19]
  reg [15:0] V1_39; // @[SWChisel.scala 164:19]
  reg [15:0] V1_40; // @[SWChisel.scala 164:19]
  reg [15:0] V1_41; // @[SWChisel.scala 164:19]
  reg [15:0] V1_42; // @[SWChisel.scala 164:19]
  reg [15:0] V1_43; // @[SWChisel.scala 164:19]
  reg [15:0] V1_44; // @[SWChisel.scala 164:19]
  reg [15:0] V1_45; // @[SWChisel.scala 164:19]
  reg [15:0] V1_46; // @[SWChisel.scala 164:19]
  reg [15:0] V1_47; // @[SWChisel.scala 164:19]
  reg [15:0] V1_48; // @[SWChisel.scala 164:19]
  reg [15:0] V1_49; // @[SWChisel.scala 164:19]
  reg [15:0] V1_50; // @[SWChisel.scala 164:19]
  reg [15:0] V1_51; // @[SWChisel.scala 164:19]
  reg [15:0] V1_52; // @[SWChisel.scala 164:19]
  reg [15:0] V1_53; // @[SWChisel.scala 164:19]
  reg [15:0] V1_54; // @[SWChisel.scala 164:19]
  reg [15:0] V1_55; // @[SWChisel.scala 164:19]
  reg [15:0] V1_56; // @[SWChisel.scala 164:19]
  reg [15:0] V1_57; // @[SWChisel.scala 164:19]
  reg [15:0] V1_58; // @[SWChisel.scala 164:19]
  reg [15:0] V1_59; // @[SWChisel.scala 164:19]
  reg [15:0] V1_60; // @[SWChisel.scala 164:19]
  reg [15:0] V2_0; // @[SWChisel.scala 166:19]
  reg [15:0] V2_1; // @[SWChisel.scala 166:19]
  reg [15:0] V2_2; // @[SWChisel.scala 166:19]
  reg [15:0] V2_3; // @[SWChisel.scala 166:19]
  reg [15:0] V2_4; // @[SWChisel.scala 166:19]
  reg [15:0] V2_5; // @[SWChisel.scala 166:19]
  reg [15:0] V2_6; // @[SWChisel.scala 166:19]
  reg [15:0] V2_7; // @[SWChisel.scala 166:19]
  reg [15:0] V2_8; // @[SWChisel.scala 166:19]
  reg [15:0] V2_9; // @[SWChisel.scala 166:19]
  reg [15:0] V2_10; // @[SWChisel.scala 166:19]
  reg [15:0] V2_11; // @[SWChisel.scala 166:19]
  reg [15:0] V2_12; // @[SWChisel.scala 166:19]
  reg [15:0] V2_13; // @[SWChisel.scala 166:19]
  reg [15:0] V2_14; // @[SWChisel.scala 166:19]
  reg [15:0] V2_15; // @[SWChisel.scala 166:19]
  reg [15:0] V2_16; // @[SWChisel.scala 166:19]
  reg [15:0] V2_17; // @[SWChisel.scala 166:19]
  reg [15:0] V2_18; // @[SWChisel.scala 166:19]
  reg [15:0] V2_19; // @[SWChisel.scala 166:19]
  reg [15:0] V2_20; // @[SWChisel.scala 166:19]
  reg [15:0] V2_21; // @[SWChisel.scala 166:19]
  reg [15:0] V2_22; // @[SWChisel.scala 166:19]
  reg [15:0] V2_23; // @[SWChisel.scala 166:19]
  reg [15:0] V2_24; // @[SWChisel.scala 166:19]
  reg [15:0] V2_25; // @[SWChisel.scala 166:19]
  reg [15:0] V2_26; // @[SWChisel.scala 166:19]
  reg [15:0] V2_27; // @[SWChisel.scala 166:19]
  reg [15:0] V2_28; // @[SWChisel.scala 166:19]
  reg [15:0] V2_29; // @[SWChisel.scala 166:19]
  reg [15:0] V2_30; // @[SWChisel.scala 166:19]
  reg [15:0] V2_31; // @[SWChisel.scala 166:19]
  reg [15:0] V2_32; // @[SWChisel.scala 166:19]
  reg [15:0] V2_33; // @[SWChisel.scala 166:19]
  reg [15:0] V2_34; // @[SWChisel.scala 166:19]
  reg [15:0] V2_35; // @[SWChisel.scala 166:19]
  reg [15:0] V2_36; // @[SWChisel.scala 166:19]
  reg [15:0] V2_37; // @[SWChisel.scala 166:19]
  reg [15:0] V2_38; // @[SWChisel.scala 166:19]
  reg [15:0] V2_39; // @[SWChisel.scala 166:19]
  reg [15:0] V2_40; // @[SWChisel.scala 166:19]
  reg [15:0] V2_41; // @[SWChisel.scala 166:19]
  reg [15:0] V2_42; // @[SWChisel.scala 166:19]
  reg [15:0] V2_43; // @[SWChisel.scala 166:19]
  reg [15:0] V2_44; // @[SWChisel.scala 166:19]
  reg [15:0] V2_45; // @[SWChisel.scala 166:19]
  reg [15:0] V2_46; // @[SWChisel.scala 166:19]
  reg [15:0] V2_47; // @[SWChisel.scala 166:19]
  reg [15:0] V2_48; // @[SWChisel.scala 166:19]
  reg [15:0] V2_49; // @[SWChisel.scala 166:19]
  reg [15:0] V2_50; // @[SWChisel.scala 166:19]
  reg [15:0] V2_51; // @[SWChisel.scala 166:19]
  reg [15:0] V2_52; // @[SWChisel.scala 166:19]
  reg [15:0] V2_53; // @[SWChisel.scala 166:19]
  reg [15:0] V2_54; // @[SWChisel.scala 166:19]
  reg [15:0] V2_55; // @[SWChisel.scala 166:19]
  reg [15:0] V2_56; // @[SWChisel.scala 166:19]
  reg [15:0] V2_57; // @[SWChisel.scala 166:19]
  reg [15:0] V2_58; // @[SWChisel.scala 166:19]
  reg [15:0] V2_59; // @[SWChisel.scala 166:19]
  reg  start_reg_0; // @[SWChisel.scala 167:26]
  reg  start_reg_1; // @[SWChisel.scala 167:26]
  reg  start_reg_2; // @[SWChisel.scala 167:26]
  reg  start_reg_3; // @[SWChisel.scala 167:26]
  reg  start_reg_4; // @[SWChisel.scala 167:26]
  reg  start_reg_5; // @[SWChisel.scala 167:26]
  reg  start_reg_6; // @[SWChisel.scala 167:26]
  reg  start_reg_7; // @[SWChisel.scala 167:26]
  reg  start_reg_8; // @[SWChisel.scala 167:26]
  reg  start_reg_9; // @[SWChisel.scala 167:26]
  reg  start_reg_10; // @[SWChisel.scala 167:26]
  reg  start_reg_11; // @[SWChisel.scala 167:26]
  reg  start_reg_12; // @[SWChisel.scala 167:26]
  reg  start_reg_13; // @[SWChisel.scala 167:26]
  reg  start_reg_14; // @[SWChisel.scala 167:26]
  reg  start_reg_15; // @[SWChisel.scala 167:26]
  reg  start_reg_16; // @[SWChisel.scala 167:26]
  reg  start_reg_17; // @[SWChisel.scala 167:26]
  reg  start_reg_18; // @[SWChisel.scala 167:26]
  reg  start_reg_19; // @[SWChisel.scala 167:26]
  reg  start_reg_20; // @[SWChisel.scala 167:26]
  reg  start_reg_21; // @[SWChisel.scala 167:26]
  reg  start_reg_22; // @[SWChisel.scala 167:26]
  reg  start_reg_23; // @[SWChisel.scala 167:26]
  reg  start_reg_24; // @[SWChisel.scala 167:26]
  reg  start_reg_25; // @[SWChisel.scala 167:26]
  reg  start_reg_26; // @[SWChisel.scala 167:26]
  reg  start_reg_27; // @[SWChisel.scala 167:26]
  reg  start_reg_28; // @[SWChisel.scala 167:26]
  reg  start_reg_29; // @[SWChisel.scala 167:26]
  reg  start_reg_30; // @[SWChisel.scala 167:26]
  reg  start_reg_31; // @[SWChisel.scala 167:26]
  reg  start_reg_32; // @[SWChisel.scala 167:26]
  reg  start_reg_33; // @[SWChisel.scala 167:26]
  reg  start_reg_34; // @[SWChisel.scala 167:26]
  reg  start_reg_35; // @[SWChisel.scala 167:26]
  reg  start_reg_36; // @[SWChisel.scala 167:26]
  reg  start_reg_37; // @[SWChisel.scala 167:26]
  reg  start_reg_38; // @[SWChisel.scala 167:26]
  reg  start_reg_39; // @[SWChisel.scala 167:26]
  reg  start_reg_40; // @[SWChisel.scala 167:26]
  reg  start_reg_41; // @[SWChisel.scala 167:26]
  reg  start_reg_42; // @[SWChisel.scala 167:26]
  reg  start_reg_43; // @[SWChisel.scala 167:26]
  reg  start_reg_44; // @[SWChisel.scala 167:26]
  reg  start_reg_45; // @[SWChisel.scala 167:26]
  reg  start_reg_46; // @[SWChisel.scala 167:26]
  reg  start_reg_47; // @[SWChisel.scala 167:26]
  reg  start_reg_48; // @[SWChisel.scala 167:26]
  reg  start_reg_49; // @[SWChisel.scala 167:26]
  reg  start_reg_50; // @[SWChisel.scala 167:26]
  reg  start_reg_51; // @[SWChisel.scala 167:26]
  reg  start_reg_52; // @[SWChisel.scala 167:26]
  reg  start_reg_53; // @[SWChisel.scala 167:26]
  reg  start_reg_54; // @[SWChisel.scala 167:26]
  reg  start_reg_55; // @[SWChisel.scala 167:26]
  reg  start_reg_56; // @[SWChisel.scala 167:26]
  reg  start_reg_57; // @[SWChisel.scala 167:26]
  reg  start_reg_58; // @[SWChisel.scala 167:26]
  reg  start_reg_59; // @[SWChisel.scala 167:26]
  wire [1:0] _GEN_181 = 9'h1 == r_count_0_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_182 = 9'h2 == r_count_0_io_out ? io_r_2_b : _GEN_181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_183 = 9'h3 == r_count_0_io_out ? io_r_3_b : _GEN_182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_184 = 9'h4 == r_count_0_io_out ? io_r_4_b : _GEN_183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_185 = 9'h5 == r_count_0_io_out ? io_r_5_b : _GEN_184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_186 = 9'h6 == r_count_0_io_out ? io_r_6_b : _GEN_185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_187 = 9'h7 == r_count_0_io_out ? io_r_7_b : _GEN_186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_188 = 9'h8 == r_count_0_io_out ? io_r_8_b : _GEN_187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_189 = 9'h9 == r_count_0_io_out ? io_r_9_b : _GEN_188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_190 = 9'ha == r_count_0_io_out ? io_r_10_b : _GEN_189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_191 = 9'hb == r_count_0_io_out ? io_r_11_b : _GEN_190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_192 = 9'hc == r_count_0_io_out ? io_r_12_b : _GEN_191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_193 = 9'hd == r_count_0_io_out ? io_r_13_b : _GEN_192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_194 = 9'he == r_count_0_io_out ? io_r_14_b : _GEN_193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_195 = 9'hf == r_count_0_io_out ? io_r_15_b : _GEN_194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_196 = 9'h10 == r_count_0_io_out ? io_r_16_b : _GEN_195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_197 = 9'h11 == r_count_0_io_out ? io_r_17_b : _GEN_196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_198 = 9'h12 == r_count_0_io_out ? io_r_18_b : _GEN_197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_199 = 9'h13 == r_count_0_io_out ? io_r_19_b : _GEN_198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_200 = 9'h14 == r_count_0_io_out ? io_r_20_b : _GEN_199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_201 = 9'h15 == r_count_0_io_out ? io_r_21_b : _GEN_200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_202 = 9'h16 == r_count_0_io_out ? io_r_22_b : _GEN_201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_203 = 9'h17 == r_count_0_io_out ? io_r_23_b : _GEN_202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_204 = 9'h18 == r_count_0_io_out ? io_r_24_b : _GEN_203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_205 = 9'h19 == r_count_0_io_out ? io_r_25_b : _GEN_204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_206 = 9'h1a == r_count_0_io_out ? io_r_26_b : _GEN_205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_207 = 9'h1b == r_count_0_io_out ? io_r_27_b : _GEN_206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_208 = 9'h1c == r_count_0_io_out ? io_r_28_b : _GEN_207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_209 = 9'h1d == r_count_0_io_out ? io_r_29_b : _GEN_208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_210 = 9'h1e == r_count_0_io_out ? io_r_30_b : _GEN_209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_211 = 9'h1f == r_count_0_io_out ? io_r_31_b : _GEN_210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_212 = 9'h20 == r_count_0_io_out ? io_r_32_b : _GEN_211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_213 = 9'h21 == r_count_0_io_out ? io_r_33_b : _GEN_212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_214 = 9'h22 == r_count_0_io_out ? io_r_34_b : _GEN_213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_215 = 9'h23 == r_count_0_io_out ? io_r_35_b : _GEN_214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_216 = 9'h24 == r_count_0_io_out ? io_r_36_b : _GEN_215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_217 = 9'h25 == r_count_0_io_out ? io_r_37_b : _GEN_216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_218 = 9'h26 == r_count_0_io_out ? io_r_38_b : _GEN_217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_219 = 9'h27 == r_count_0_io_out ? io_r_39_b : _GEN_218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_220 = 9'h28 == r_count_0_io_out ? io_r_40_b : _GEN_219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_221 = 9'h29 == r_count_0_io_out ? io_r_41_b : _GEN_220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_222 = 9'h2a == r_count_0_io_out ? io_r_42_b : _GEN_221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_223 = 9'h2b == r_count_0_io_out ? io_r_43_b : _GEN_222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_224 = 9'h2c == r_count_0_io_out ? io_r_44_b : _GEN_223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_225 = 9'h2d == r_count_0_io_out ? io_r_45_b : _GEN_224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_226 = 9'h2e == r_count_0_io_out ? io_r_46_b : _GEN_225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_227 = 9'h2f == r_count_0_io_out ? io_r_47_b : _GEN_226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_228 = 9'h30 == r_count_0_io_out ? io_r_48_b : _GEN_227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_229 = 9'h31 == r_count_0_io_out ? io_r_49_b : _GEN_228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_230 = 9'h32 == r_count_0_io_out ? io_r_50_b : _GEN_229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_231 = 9'h33 == r_count_0_io_out ? io_r_51_b : _GEN_230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_232 = 9'h34 == r_count_0_io_out ? io_r_52_b : _GEN_231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_233 = 9'h35 == r_count_0_io_out ? io_r_53_b : _GEN_232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_234 = 9'h36 == r_count_0_io_out ? io_r_54_b : _GEN_233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_235 = 9'h37 == r_count_0_io_out ? io_r_55_b : _GEN_234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_236 = 9'h38 == r_count_0_io_out ? io_r_56_b : _GEN_235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_237 = 9'h39 == r_count_0_io_out ? io_r_57_b : _GEN_236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_238 = 9'h3a == r_count_0_io_out ? io_r_58_b : _GEN_237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_239 = 9'h3b == r_count_0_io_out ? io_r_59_b : _GEN_238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_240 = 9'h3c == r_count_0_io_out ? io_r_60_b : _GEN_239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_241 = 9'h3d == r_count_0_io_out ? io_r_61_b : _GEN_240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_242 = 9'h3e == r_count_0_io_out ? io_r_62_b : _GEN_241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_243 = 9'h3f == r_count_0_io_out ? io_r_63_b : _GEN_242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_244 = 9'h40 == r_count_0_io_out ? io_r_64_b : _GEN_243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_245 = 9'h41 == r_count_0_io_out ? io_r_65_b : _GEN_244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_246 = 9'h42 == r_count_0_io_out ? io_r_66_b : _GEN_245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_247 = 9'h43 == r_count_0_io_out ? io_r_67_b : _GEN_246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_248 = 9'h44 == r_count_0_io_out ? io_r_68_b : _GEN_247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_249 = 9'h45 == r_count_0_io_out ? io_r_69_b : _GEN_248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_250 = 9'h46 == r_count_0_io_out ? io_r_70_b : _GEN_249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_251 = 9'h47 == r_count_0_io_out ? io_r_71_b : _GEN_250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_252 = 9'h48 == r_count_0_io_out ? io_r_72_b : _GEN_251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_253 = 9'h49 == r_count_0_io_out ? io_r_73_b : _GEN_252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_254 = 9'h4a == r_count_0_io_out ? io_r_74_b : _GEN_253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_255 = 9'h4b == r_count_0_io_out ? io_r_75_b : _GEN_254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_256 = 9'h4c == r_count_0_io_out ? io_r_76_b : _GEN_255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_257 = 9'h4d == r_count_0_io_out ? io_r_77_b : _GEN_256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_258 = 9'h4e == r_count_0_io_out ? io_r_78_b : _GEN_257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_259 = 9'h4f == r_count_0_io_out ? io_r_79_b : _GEN_258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_260 = 9'h50 == r_count_0_io_out ? io_r_80_b : _GEN_259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_261 = 9'h51 == r_count_0_io_out ? io_r_81_b : _GEN_260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_262 = 9'h52 == r_count_0_io_out ? io_r_82_b : _GEN_261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_263 = 9'h53 == r_count_0_io_out ? io_r_83_b : _GEN_262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_264 = 9'h54 == r_count_0_io_out ? io_r_84_b : _GEN_263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_265 = 9'h55 == r_count_0_io_out ? io_r_85_b : _GEN_264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_266 = 9'h56 == r_count_0_io_out ? io_r_86_b : _GEN_265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_267 = 9'h57 == r_count_0_io_out ? io_r_87_b : _GEN_266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_268 = 9'h58 == r_count_0_io_out ? io_r_88_b : _GEN_267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_269 = 9'h59 == r_count_0_io_out ? io_r_89_b : _GEN_268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_270 = 9'h5a == r_count_0_io_out ? io_r_90_b : _GEN_269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_271 = 9'h5b == r_count_0_io_out ? io_r_91_b : _GEN_270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_272 = 9'h5c == r_count_0_io_out ? io_r_92_b : _GEN_271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_273 = 9'h5d == r_count_0_io_out ? io_r_93_b : _GEN_272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_274 = 9'h5e == r_count_0_io_out ? io_r_94_b : _GEN_273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_275 = 9'h5f == r_count_0_io_out ? io_r_95_b : _GEN_274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_276 = 9'h60 == r_count_0_io_out ? io_r_96_b : _GEN_275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_277 = 9'h61 == r_count_0_io_out ? io_r_97_b : _GEN_276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_278 = 9'h62 == r_count_0_io_out ? io_r_98_b : _GEN_277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_279 = 9'h63 == r_count_0_io_out ? io_r_99_b : _GEN_278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_280 = 9'h64 == r_count_0_io_out ? io_r_100_b : _GEN_279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_281 = 9'h65 == r_count_0_io_out ? io_r_101_b : _GEN_280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_282 = 9'h66 == r_count_0_io_out ? io_r_102_b : _GEN_281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_283 = 9'h67 == r_count_0_io_out ? io_r_103_b : _GEN_282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_284 = 9'h68 == r_count_0_io_out ? io_r_104_b : _GEN_283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_285 = 9'h69 == r_count_0_io_out ? io_r_105_b : _GEN_284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_286 = 9'h6a == r_count_0_io_out ? io_r_106_b : _GEN_285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_287 = 9'h6b == r_count_0_io_out ? io_r_107_b : _GEN_286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_288 = 9'h6c == r_count_0_io_out ? io_r_108_b : _GEN_287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_289 = 9'h6d == r_count_0_io_out ? io_r_109_b : _GEN_288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_290 = 9'h6e == r_count_0_io_out ? io_r_110_b : _GEN_289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_291 = 9'h6f == r_count_0_io_out ? io_r_111_b : _GEN_290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_292 = 9'h70 == r_count_0_io_out ? io_r_112_b : _GEN_291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_293 = 9'h71 == r_count_0_io_out ? io_r_113_b : _GEN_292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_294 = 9'h72 == r_count_0_io_out ? io_r_114_b : _GEN_293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_295 = 9'h73 == r_count_0_io_out ? io_r_115_b : _GEN_294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_296 = 9'h74 == r_count_0_io_out ? io_r_116_b : _GEN_295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_297 = 9'h75 == r_count_0_io_out ? io_r_117_b : _GEN_296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_298 = 9'h76 == r_count_0_io_out ? io_r_118_b : _GEN_297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_299 = 9'h77 == r_count_0_io_out ? io_r_119_b : _GEN_298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_300 = 9'h78 == r_count_0_io_out ? io_r_120_b : _GEN_299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_301 = 9'h79 == r_count_0_io_out ? io_r_121_b : _GEN_300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_302 = 9'h7a == r_count_0_io_out ? io_r_122_b : _GEN_301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_303 = 9'h7b == r_count_0_io_out ? io_r_123_b : _GEN_302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_304 = 9'h7c == r_count_0_io_out ? io_r_124_b : _GEN_303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_305 = 9'h7d == r_count_0_io_out ? io_r_125_b : _GEN_304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_306 = 9'h7e == r_count_0_io_out ? io_r_126_b : _GEN_305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_307 = 9'h7f == r_count_0_io_out ? io_r_127_b : _GEN_306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_308 = 9'h80 == r_count_0_io_out ? io_r_128_b : _GEN_307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_309 = 9'h81 == r_count_0_io_out ? io_r_129_b : _GEN_308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_310 = 9'h82 == r_count_0_io_out ? io_r_130_b : _GEN_309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_311 = 9'h83 == r_count_0_io_out ? io_r_131_b : _GEN_310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_312 = 9'h84 == r_count_0_io_out ? io_r_132_b : _GEN_311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_313 = 9'h85 == r_count_0_io_out ? io_r_133_b : _GEN_312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_314 = 9'h86 == r_count_0_io_out ? io_r_134_b : _GEN_313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_315 = 9'h87 == r_count_0_io_out ? io_r_135_b : _GEN_314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_316 = 9'h88 == r_count_0_io_out ? io_r_136_b : _GEN_315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_317 = 9'h89 == r_count_0_io_out ? io_r_137_b : _GEN_316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_318 = 9'h8a == r_count_0_io_out ? io_r_138_b : _GEN_317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_319 = 9'h8b == r_count_0_io_out ? io_r_139_b : _GEN_318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_320 = 9'h8c == r_count_0_io_out ? io_r_140_b : _GEN_319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_321 = 9'h8d == r_count_0_io_out ? io_r_141_b : _GEN_320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_322 = 9'h8e == r_count_0_io_out ? io_r_142_b : _GEN_321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_323 = 9'h8f == r_count_0_io_out ? io_r_143_b : _GEN_322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_324 = 9'h90 == r_count_0_io_out ? io_r_144_b : _GEN_323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_325 = 9'h91 == r_count_0_io_out ? io_r_145_b : _GEN_324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_326 = 9'h92 == r_count_0_io_out ? io_r_146_b : _GEN_325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_327 = 9'h93 == r_count_0_io_out ? io_r_147_b : _GEN_326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_328 = 9'h94 == r_count_0_io_out ? io_r_148_b : _GEN_327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_329 = 9'h95 == r_count_0_io_out ? io_r_149_b : _GEN_328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_330 = 9'h96 == r_count_0_io_out ? io_r_150_b : _GEN_329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_331 = 9'h97 == r_count_0_io_out ? io_r_151_b : _GEN_330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_332 = 9'h98 == r_count_0_io_out ? io_r_152_b : _GEN_331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_333 = 9'h99 == r_count_0_io_out ? io_r_153_b : _GEN_332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_334 = 9'h9a == r_count_0_io_out ? io_r_154_b : _GEN_333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_335 = 9'h9b == r_count_0_io_out ? io_r_155_b : _GEN_334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_336 = 9'h9c == r_count_0_io_out ? io_r_156_b : _GEN_335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_337 = 9'h9d == r_count_0_io_out ? io_r_157_b : _GEN_336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_338 = 9'h9e == r_count_0_io_out ? io_r_158_b : _GEN_337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_339 = 9'h9f == r_count_0_io_out ? io_r_159_b : _GEN_338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_340 = 9'ha0 == r_count_0_io_out ? io_r_160_b : _GEN_339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_341 = 9'ha1 == r_count_0_io_out ? io_r_161_b : _GEN_340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_342 = 9'ha2 == r_count_0_io_out ? io_r_162_b : _GEN_341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_343 = 9'ha3 == r_count_0_io_out ? io_r_163_b : _GEN_342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_344 = 9'ha4 == r_count_0_io_out ? io_r_164_b : _GEN_343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_345 = 9'ha5 == r_count_0_io_out ? io_r_165_b : _GEN_344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_346 = 9'ha6 == r_count_0_io_out ? io_r_166_b : _GEN_345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_347 = 9'ha7 == r_count_0_io_out ? io_r_167_b : _GEN_346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_348 = 9'ha8 == r_count_0_io_out ? io_r_168_b : _GEN_347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_349 = 9'ha9 == r_count_0_io_out ? io_r_169_b : _GEN_348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_350 = 9'haa == r_count_0_io_out ? io_r_170_b : _GEN_349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_351 = 9'hab == r_count_0_io_out ? io_r_171_b : _GEN_350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_352 = 9'hac == r_count_0_io_out ? io_r_172_b : _GEN_351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_353 = 9'had == r_count_0_io_out ? io_r_173_b : _GEN_352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_354 = 9'hae == r_count_0_io_out ? io_r_174_b : _GEN_353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_355 = 9'haf == r_count_0_io_out ? io_r_175_b : _GEN_354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_356 = 9'hb0 == r_count_0_io_out ? io_r_176_b : _GEN_355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_357 = 9'hb1 == r_count_0_io_out ? io_r_177_b : _GEN_356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_358 = 9'hb2 == r_count_0_io_out ? io_r_178_b : _GEN_357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_359 = 9'hb3 == r_count_0_io_out ? io_r_179_b : _GEN_358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_360 = 9'hb4 == r_count_0_io_out ? io_r_180_b : _GEN_359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_361 = 9'hb5 == r_count_0_io_out ? io_r_181_b : _GEN_360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_362 = 9'hb6 == r_count_0_io_out ? io_r_182_b : _GEN_361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_363 = 9'hb7 == r_count_0_io_out ? io_r_183_b : _GEN_362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_364 = 9'hb8 == r_count_0_io_out ? io_r_184_b : _GEN_363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_365 = 9'hb9 == r_count_0_io_out ? io_r_185_b : _GEN_364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_366 = 9'hba == r_count_0_io_out ? io_r_186_b : _GEN_365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_367 = 9'hbb == r_count_0_io_out ? io_r_187_b : _GEN_366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_368 = 9'hbc == r_count_0_io_out ? io_r_188_b : _GEN_367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_369 = 9'hbd == r_count_0_io_out ? io_r_189_b : _GEN_368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_370 = 9'hbe == r_count_0_io_out ? io_r_190_b : _GEN_369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_371 = 9'hbf == r_count_0_io_out ? io_r_191_b : _GEN_370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_372 = 9'hc0 == r_count_0_io_out ? io_r_192_b : _GEN_371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_373 = 9'hc1 == r_count_0_io_out ? io_r_193_b : _GEN_372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_374 = 9'hc2 == r_count_0_io_out ? io_r_194_b : _GEN_373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_375 = 9'hc3 == r_count_0_io_out ? io_r_195_b : _GEN_374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_376 = 9'hc4 == r_count_0_io_out ? io_r_196_b : _GEN_375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_377 = 9'hc5 == r_count_0_io_out ? io_r_197_b : _GEN_376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_378 = 9'hc6 == r_count_0_io_out ? io_r_198_b : _GEN_377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_379 = 9'hc7 == r_count_0_io_out ? io_r_199_b : _GEN_378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_380 = 9'hc8 == r_count_0_io_out ? io_r_200_b : _GEN_379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_381 = 9'hc9 == r_count_0_io_out ? io_r_201_b : _GEN_380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_382 = 9'hca == r_count_0_io_out ? io_r_202_b : _GEN_381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_383 = 9'hcb == r_count_0_io_out ? io_r_203_b : _GEN_382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_384 = 9'hcc == r_count_0_io_out ? io_r_204_b : _GEN_383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_385 = 9'hcd == r_count_0_io_out ? io_r_205_b : _GEN_384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_386 = 9'hce == r_count_0_io_out ? io_r_206_b : _GEN_385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_387 = 9'hcf == r_count_0_io_out ? io_r_207_b : _GEN_386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_388 = 9'hd0 == r_count_0_io_out ? io_r_208_b : _GEN_387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_389 = 9'hd1 == r_count_0_io_out ? io_r_209_b : _GEN_388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_390 = 9'hd2 == r_count_0_io_out ? io_r_210_b : _GEN_389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_391 = 9'hd3 == r_count_0_io_out ? io_r_211_b : _GEN_390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_392 = 9'hd4 == r_count_0_io_out ? io_r_212_b : _GEN_391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_393 = 9'hd5 == r_count_0_io_out ? io_r_213_b : _GEN_392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_394 = 9'hd6 == r_count_0_io_out ? io_r_214_b : _GEN_393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_395 = 9'hd7 == r_count_0_io_out ? io_r_215_b : _GEN_394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_396 = 9'hd8 == r_count_0_io_out ? io_r_216_b : _GEN_395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_397 = 9'hd9 == r_count_0_io_out ? io_r_217_b : _GEN_396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_398 = 9'hda == r_count_0_io_out ? io_r_218_b : _GEN_397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_399 = 9'hdb == r_count_0_io_out ? io_r_219_b : _GEN_398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_400 = 9'hdc == r_count_0_io_out ? io_r_220_b : _GEN_399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_401 = 9'hdd == r_count_0_io_out ? io_r_221_b : _GEN_400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_402 = 9'hde == r_count_0_io_out ? io_r_222_b : _GEN_401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_403 = 9'hdf == r_count_0_io_out ? io_r_223_b : _GEN_402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_404 = 9'he0 == r_count_0_io_out ? io_r_224_b : _GEN_403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_405 = 9'he1 == r_count_0_io_out ? io_r_225_b : _GEN_404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_406 = 9'he2 == r_count_0_io_out ? io_r_226_b : _GEN_405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_407 = 9'he3 == r_count_0_io_out ? io_r_227_b : _GEN_406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_408 = 9'he4 == r_count_0_io_out ? io_r_228_b : _GEN_407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_409 = 9'he5 == r_count_0_io_out ? io_r_229_b : _GEN_408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_410 = 9'he6 == r_count_0_io_out ? io_r_230_b : _GEN_409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_411 = 9'he7 == r_count_0_io_out ? io_r_231_b : _GEN_410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_412 = 9'he8 == r_count_0_io_out ? io_r_232_b : _GEN_411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_413 = 9'he9 == r_count_0_io_out ? io_r_233_b : _GEN_412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_414 = 9'hea == r_count_0_io_out ? io_r_234_b : _GEN_413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_415 = 9'heb == r_count_0_io_out ? io_r_235_b : _GEN_414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_416 = 9'hec == r_count_0_io_out ? io_r_236_b : _GEN_415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_417 = 9'hed == r_count_0_io_out ? io_r_237_b : _GEN_416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_418 = 9'hee == r_count_0_io_out ? io_r_238_b : _GEN_417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_419 = 9'hef == r_count_0_io_out ? io_r_239_b : _GEN_418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_420 = 9'hf0 == r_count_0_io_out ? io_r_240_b : _GEN_419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_421 = 9'hf1 == r_count_0_io_out ? io_r_241_b : _GEN_420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_422 = 9'hf2 == r_count_0_io_out ? io_r_242_b : _GEN_421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_423 = 9'hf3 == r_count_0_io_out ? io_r_243_b : _GEN_422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_424 = 9'hf4 == r_count_0_io_out ? io_r_244_b : _GEN_423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_425 = 9'hf5 == r_count_0_io_out ? io_r_245_b : _GEN_424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_426 = 9'hf6 == r_count_0_io_out ? io_r_246_b : _GEN_425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_427 = 9'hf7 == r_count_0_io_out ? io_r_247_b : _GEN_426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_428 = 9'hf8 == r_count_0_io_out ? io_r_248_b : _GEN_427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_429 = 9'hf9 == r_count_0_io_out ? io_r_249_b : _GEN_428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_430 = 9'hfa == r_count_0_io_out ? io_r_250_b : _GEN_429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_431 = 9'hfb == r_count_0_io_out ? io_r_251_b : _GEN_430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_432 = 9'hfc == r_count_0_io_out ? io_r_252_b : _GEN_431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_433 = 9'hfd == r_count_0_io_out ? io_r_253_b : _GEN_432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_434 = 9'hfe == r_count_0_io_out ? io_r_254_b : _GEN_433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_435 = 9'hff == r_count_0_io_out ? io_r_255_b : _GEN_434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_436 = 9'h100 == r_count_0_io_out ? io_r_256_b : _GEN_435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_437 = 9'h101 == r_count_0_io_out ? io_r_257_b : _GEN_436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_438 = 9'h102 == r_count_0_io_out ? io_r_258_b : _GEN_437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_439 = 9'h103 == r_count_0_io_out ? io_r_259_b : _GEN_438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_440 = 9'h104 == r_count_0_io_out ? io_r_260_b : _GEN_439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_441 = 9'h105 == r_count_0_io_out ? io_r_261_b : _GEN_440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_442 = 9'h106 == r_count_0_io_out ? io_r_262_b : _GEN_441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_443 = 9'h107 == r_count_0_io_out ? io_r_263_b : _GEN_442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_444 = 9'h108 == r_count_0_io_out ? io_r_264_b : _GEN_443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_445 = 9'h109 == r_count_0_io_out ? io_r_265_b : _GEN_444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_446 = 9'h10a == r_count_0_io_out ? io_r_266_b : _GEN_445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_447 = 9'h10b == r_count_0_io_out ? io_r_267_b : _GEN_446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_448 = 9'h10c == r_count_0_io_out ? io_r_268_b : _GEN_447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_449 = 9'h10d == r_count_0_io_out ? io_r_269_b : _GEN_448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_450 = 9'h10e == r_count_0_io_out ? io_r_270_b : _GEN_449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_451 = 9'h10f == r_count_0_io_out ? io_r_271_b : _GEN_450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_452 = 9'h110 == r_count_0_io_out ? io_r_272_b : _GEN_451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_453 = 9'h111 == r_count_0_io_out ? io_r_273_b : _GEN_452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_454 = 9'h112 == r_count_0_io_out ? io_r_274_b : _GEN_453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_455 = 9'h113 == r_count_0_io_out ? io_r_275_b : _GEN_454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_456 = 9'h114 == r_count_0_io_out ? io_r_276_b : _GEN_455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_457 = 9'h115 == r_count_0_io_out ? io_r_277_b : _GEN_456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_458 = 9'h116 == r_count_0_io_out ? io_r_278_b : _GEN_457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_459 = 9'h117 == r_count_0_io_out ? io_r_279_b : _GEN_458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_460 = 9'h118 == r_count_0_io_out ? io_r_280_b : _GEN_459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_461 = 9'h119 == r_count_0_io_out ? io_r_281_b : _GEN_460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_462 = 9'h11a == r_count_0_io_out ? io_r_282_b : _GEN_461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_463 = 9'h11b == r_count_0_io_out ? io_r_283_b : _GEN_462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_464 = 9'h11c == r_count_0_io_out ? io_r_284_b : _GEN_463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_465 = 9'h11d == r_count_0_io_out ? io_r_285_b : _GEN_464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_466 = 9'h11e == r_count_0_io_out ? io_r_286_b : _GEN_465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_467 = 9'h11f == r_count_0_io_out ? io_r_287_b : _GEN_466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_468 = 9'h120 == r_count_0_io_out ? io_r_288_b : _GEN_467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_469 = 9'h121 == r_count_0_io_out ? io_r_289_b : _GEN_468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_470 = 9'h122 == r_count_0_io_out ? io_r_290_b : _GEN_469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_471 = 9'h123 == r_count_0_io_out ? io_r_291_b : _GEN_470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_472 = 9'h124 == r_count_0_io_out ? io_r_292_b : _GEN_471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_473 = 9'h125 == r_count_0_io_out ? io_r_293_b : _GEN_472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_474 = 9'h126 == r_count_0_io_out ? io_r_294_b : _GEN_473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_475 = 9'h127 == r_count_0_io_out ? io_r_295_b : _GEN_474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_476 = 9'h128 == r_count_0_io_out ? io_r_296_b : _GEN_475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_477 = 9'h129 == r_count_0_io_out ? io_r_297_b : _GEN_476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_478 = 9'h12a == r_count_0_io_out ? io_r_298_b : _GEN_477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_479 = 9'h12b == r_count_0_io_out ? io_r_299_b : _GEN_478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_480 = 9'h12c == r_count_0_io_out ? io_r_300_b : _GEN_479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_481 = 9'h12d == r_count_0_io_out ? io_r_301_b : _GEN_480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_482 = 9'h12e == r_count_0_io_out ? io_r_302_b : _GEN_481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_483 = 9'h12f == r_count_0_io_out ? io_r_303_b : _GEN_482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_484 = 9'h130 == r_count_0_io_out ? io_r_304_b : _GEN_483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_485 = 9'h131 == r_count_0_io_out ? io_r_305_b : _GEN_484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_486 = 9'h132 == r_count_0_io_out ? io_r_306_b : _GEN_485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_487 = 9'h133 == r_count_0_io_out ? io_r_307_b : _GEN_486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_488 = 9'h134 == r_count_0_io_out ? io_r_308_b : _GEN_487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_489 = 9'h135 == r_count_0_io_out ? io_r_309_b : _GEN_488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_490 = 9'h136 == r_count_0_io_out ? io_r_310_b : _GEN_489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_491 = 9'h137 == r_count_0_io_out ? io_r_311_b : _GEN_490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_492 = 9'h138 == r_count_0_io_out ? io_r_312_b : _GEN_491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_493 = 9'h139 == r_count_0_io_out ? io_r_313_b : _GEN_492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_494 = 9'h13a == r_count_0_io_out ? io_r_314_b : _GEN_493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_495 = 9'h13b == r_count_0_io_out ? io_r_315_b : _GEN_494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_496 = 9'h13c == r_count_0_io_out ? io_r_316_b : _GEN_495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_497 = 9'h13d == r_count_0_io_out ? io_r_317_b : _GEN_496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_498 = 9'h13e == r_count_0_io_out ? io_r_318_b : _GEN_497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_499 = 9'h13f == r_count_0_io_out ? io_r_319_b : _GEN_498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_500 = 9'h140 == r_count_0_io_out ? io_r_320_b : _GEN_499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_501 = 9'h141 == r_count_0_io_out ? io_r_321_b : _GEN_500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_502 = 9'h142 == r_count_0_io_out ? io_r_322_b : _GEN_501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_503 = 9'h143 == r_count_0_io_out ? io_r_323_b : _GEN_502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_504 = 9'h144 == r_count_0_io_out ? io_r_324_b : _GEN_503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_505 = 9'h145 == r_count_0_io_out ? io_r_325_b : _GEN_504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_506 = 9'h146 == r_count_0_io_out ? io_r_326_b : _GEN_505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_507 = 9'h147 == r_count_0_io_out ? io_r_327_b : _GEN_506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_508 = 9'h148 == r_count_0_io_out ? io_r_328_b : _GEN_507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_509 = 9'h149 == r_count_0_io_out ? io_r_329_b : _GEN_508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_510 = 9'h14a == r_count_0_io_out ? io_r_330_b : _GEN_509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_511 = 9'h14b == r_count_0_io_out ? io_r_331_b : _GEN_510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_512 = 9'h14c == r_count_0_io_out ? io_r_332_b : _GEN_511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_513 = 9'h14d == r_count_0_io_out ? io_r_333_b : _GEN_512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_514 = 9'h14e == r_count_0_io_out ? io_r_334_b : _GEN_513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_515 = 9'h14f == r_count_0_io_out ? io_r_335_b : _GEN_514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_516 = 9'h150 == r_count_0_io_out ? io_r_336_b : _GEN_515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_517 = 9'h151 == r_count_0_io_out ? io_r_337_b : _GEN_516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_518 = 9'h152 == r_count_0_io_out ? io_r_338_b : _GEN_517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_519 = 9'h153 == r_count_0_io_out ? io_r_339_b : _GEN_518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_520 = 9'h154 == r_count_0_io_out ? io_r_340_b : _GEN_519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_521 = 9'h155 == r_count_0_io_out ? io_r_341_b : _GEN_520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_522 = 9'h156 == r_count_0_io_out ? io_r_342_b : _GEN_521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_523 = 9'h157 == r_count_0_io_out ? io_r_343_b : _GEN_522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_524 = 9'h158 == r_count_0_io_out ? io_r_344_b : _GEN_523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_525 = 9'h159 == r_count_0_io_out ? io_r_345_b : _GEN_524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_526 = 9'h15a == r_count_0_io_out ? io_r_346_b : _GEN_525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_527 = 9'h15b == r_count_0_io_out ? io_r_347_b : _GEN_526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_528 = 9'h15c == r_count_0_io_out ? io_r_348_b : _GEN_527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_529 = 9'h15d == r_count_0_io_out ? io_r_349_b : _GEN_528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_530 = 9'h15e == r_count_0_io_out ? io_r_350_b : _GEN_529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_531 = 9'h15f == r_count_0_io_out ? io_r_351_b : _GEN_530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_532 = 9'h160 == r_count_0_io_out ? io_r_352_b : _GEN_531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_533 = 9'h161 == r_count_0_io_out ? io_r_353_b : _GEN_532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_534 = 9'h162 == r_count_0_io_out ? io_r_354_b : _GEN_533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_535 = 9'h163 == r_count_0_io_out ? io_r_355_b : _GEN_534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_536 = 9'h164 == r_count_0_io_out ? io_r_356_b : _GEN_535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_537 = 9'h165 == r_count_0_io_out ? io_r_357_b : _GEN_536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_538 = 9'h166 == r_count_0_io_out ? io_r_358_b : _GEN_537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_539 = 9'h167 == r_count_0_io_out ? io_r_359_b : _GEN_538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_540 = 9'h168 == r_count_0_io_out ? io_r_360_b : _GEN_539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_541 = 9'h169 == r_count_0_io_out ? io_r_361_b : _GEN_540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_542 = 9'h16a == r_count_0_io_out ? io_r_362_b : _GEN_541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_543 = 9'h16b == r_count_0_io_out ? io_r_363_b : _GEN_542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_544 = 9'h16c == r_count_0_io_out ? io_r_364_b : _GEN_543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_545 = 9'h16d == r_count_0_io_out ? io_r_365_b : _GEN_544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_546 = 9'h16e == r_count_0_io_out ? io_r_366_b : _GEN_545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_547 = 9'h16f == r_count_0_io_out ? io_r_367_b : _GEN_546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_548 = 9'h170 == r_count_0_io_out ? io_r_368_b : _GEN_547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_549 = 9'h171 == r_count_0_io_out ? io_r_369_b : _GEN_548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_550 = 9'h172 == r_count_0_io_out ? io_r_370_b : _GEN_549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_551 = 9'h173 == r_count_0_io_out ? io_r_371_b : _GEN_550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_552 = 9'h174 == r_count_0_io_out ? io_r_372_b : _GEN_551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_553 = 9'h175 == r_count_0_io_out ? io_r_373_b : _GEN_552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_554 = 9'h176 == r_count_0_io_out ? io_r_374_b : _GEN_553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_555 = 9'h177 == r_count_0_io_out ? io_r_375_b : _GEN_554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_556 = 9'h178 == r_count_0_io_out ? io_r_376_b : _GEN_555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_557 = 9'h179 == r_count_0_io_out ? io_r_377_b : _GEN_556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_558 = 9'h17a == r_count_0_io_out ? io_r_378_b : _GEN_557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_559 = 9'h17b == r_count_0_io_out ? io_r_379_b : _GEN_558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_560 = 9'h17c == r_count_0_io_out ? io_r_380_b : _GEN_559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_561 = 9'h17d == r_count_0_io_out ? io_r_381_b : _GEN_560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_562 = 9'h17e == r_count_0_io_out ? io_r_382_b : _GEN_561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_563 = 9'h17f == r_count_0_io_out ? io_r_383_b : _GEN_562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_564 = 9'h180 == r_count_0_io_out ? io_r_384_b : _GEN_563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_565 = 9'h181 == r_count_0_io_out ? io_r_385_b : _GEN_564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_566 = 9'h182 == r_count_0_io_out ? io_r_386_b : _GEN_565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_567 = 9'h183 == r_count_0_io_out ? io_r_387_b : _GEN_566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_568 = 9'h184 == r_count_0_io_out ? io_r_388_b : _GEN_567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_569 = 9'h185 == r_count_0_io_out ? io_r_389_b : _GEN_568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_570 = 9'h186 == r_count_0_io_out ? io_r_390_b : _GEN_569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_571 = 9'h187 == r_count_0_io_out ? io_r_391_b : _GEN_570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_572 = 9'h188 == r_count_0_io_out ? io_r_392_b : _GEN_571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_573 = 9'h189 == r_count_0_io_out ? io_r_393_b : _GEN_572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_574 = 9'h18a == r_count_0_io_out ? io_r_394_b : _GEN_573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_575 = 9'h18b == r_count_0_io_out ? io_r_395_b : _GEN_574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_576 = 9'h18c == r_count_0_io_out ? io_r_396_b : _GEN_575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_577 = 9'h18d == r_count_0_io_out ? io_r_397_b : _GEN_576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_578 = 9'h18e == r_count_0_io_out ? io_r_398_b : _GEN_577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_581 = 9'h1 == r_count_1_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_582 = 9'h2 == r_count_1_io_out ? io_r_2_b : _GEN_581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_583 = 9'h3 == r_count_1_io_out ? io_r_3_b : _GEN_582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_584 = 9'h4 == r_count_1_io_out ? io_r_4_b : _GEN_583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_585 = 9'h5 == r_count_1_io_out ? io_r_5_b : _GEN_584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_586 = 9'h6 == r_count_1_io_out ? io_r_6_b : _GEN_585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_587 = 9'h7 == r_count_1_io_out ? io_r_7_b : _GEN_586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_588 = 9'h8 == r_count_1_io_out ? io_r_8_b : _GEN_587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_589 = 9'h9 == r_count_1_io_out ? io_r_9_b : _GEN_588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_590 = 9'ha == r_count_1_io_out ? io_r_10_b : _GEN_589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_591 = 9'hb == r_count_1_io_out ? io_r_11_b : _GEN_590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_592 = 9'hc == r_count_1_io_out ? io_r_12_b : _GEN_591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_593 = 9'hd == r_count_1_io_out ? io_r_13_b : _GEN_592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_594 = 9'he == r_count_1_io_out ? io_r_14_b : _GEN_593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_595 = 9'hf == r_count_1_io_out ? io_r_15_b : _GEN_594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_596 = 9'h10 == r_count_1_io_out ? io_r_16_b : _GEN_595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_597 = 9'h11 == r_count_1_io_out ? io_r_17_b : _GEN_596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_598 = 9'h12 == r_count_1_io_out ? io_r_18_b : _GEN_597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_599 = 9'h13 == r_count_1_io_out ? io_r_19_b : _GEN_598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_600 = 9'h14 == r_count_1_io_out ? io_r_20_b : _GEN_599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_601 = 9'h15 == r_count_1_io_out ? io_r_21_b : _GEN_600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_602 = 9'h16 == r_count_1_io_out ? io_r_22_b : _GEN_601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_603 = 9'h17 == r_count_1_io_out ? io_r_23_b : _GEN_602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_604 = 9'h18 == r_count_1_io_out ? io_r_24_b : _GEN_603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_605 = 9'h19 == r_count_1_io_out ? io_r_25_b : _GEN_604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_606 = 9'h1a == r_count_1_io_out ? io_r_26_b : _GEN_605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_607 = 9'h1b == r_count_1_io_out ? io_r_27_b : _GEN_606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_608 = 9'h1c == r_count_1_io_out ? io_r_28_b : _GEN_607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_609 = 9'h1d == r_count_1_io_out ? io_r_29_b : _GEN_608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_610 = 9'h1e == r_count_1_io_out ? io_r_30_b : _GEN_609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_611 = 9'h1f == r_count_1_io_out ? io_r_31_b : _GEN_610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_612 = 9'h20 == r_count_1_io_out ? io_r_32_b : _GEN_611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_613 = 9'h21 == r_count_1_io_out ? io_r_33_b : _GEN_612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_614 = 9'h22 == r_count_1_io_out ? io_r_34_b : _GEN_613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_615 = 9'h23 == r_count_1_io_out ? io_r_35_b : _GEN_614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_616 = 9'h24 == r_count_1_io_out ? io_r_36_b : _GEN_615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_617 = 9'h25 == r_count_1_io_out ? io_r_37_b : _GEN_616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_618 = 9'h26 == r_count_1_io_out ? io_r_38_b : _GEN_617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_619 = 9'h27 == r_count_1_io_out ? io_r_39_b : _GEN_618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_620 = 9'h28 == r_count_1_io_out ? io_r_40_b : _GEN_619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_621 = 9'h29 == r_count_1_io_out ? io_r_41_b : _GEN_620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_622 = 9'h2a == r_count_1_io_out ? io_r_42_b : _GEN_621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_623 = 9'h2b == r_count_1_io_out ? io_r_43_b : _GEN_622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_624 = 9'h2c == r_count_1_io_out ? io_r_44_b : _GEN_623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_625 = 9'h2d == r_count_1_io_out ? io_r_45_b : _GEN_624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_626 = 9'h2e == r_count_1_io_out ? io_r_46_b : _GEN_625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_627 = 9'h2f == r_count_1_io_out ? io_r_47_b : _GEN_626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_628 = 9'h30 == r_count_1_io_out ? io_r_48_b : _GEN_627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_629 = 9'h31 == r_count_1_io_out ? io_r_49_b : _GEN_628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_630 = 9'h32 == r_count_1_io_out ? io_r_50_b : _GEN_629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_631 = 9'h33 == r_count_1_io_out ? io_r_51_b : _GEN_630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_632 = 9'h34 == r_count_1_io_out ? io_r_52_b : _GEN_631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_633 = 9'h35 == r_count_1_io_out ? io_r_53_b : _GEN_632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_634 = 9'h36 == r_count_1_io_out ? io_r_54_b : _GEN_633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_635 = 9'h37 == r_count_1_io_out ? io_r_55_b : _GEN_634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_636 = 9'h38 == r_count_1_io_out ? io_r_56_b : _GEN_635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_637 = 9'h39 == r_count_1_io_out ? io_r_57_b : _GEN_636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_638 = 9'h3a == r_count_1_io_out ? io_r_58_b : _GEN_637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_639 = 9'h3b == r_count_1_io_out ? io_r_59_b : _GEN_638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_640 = 9'h3c == r_count_1_io_out ? io_r_60_b : _GEN_639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_641 = 9'h3d == r_count_1_io_out ? io_r_61_b : _GEN_640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_642 = 9'h3e == r_count_1_io_out ? io_r_62_b : _GEN_641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_643 = 9'h3f == r_count_1_io_out ? io_r_63_b : _GEN_642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_644 = 9'h40 == r_count_1_io_out ? io_r_64_b : _GEN_643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_645 = 9'h41 == r_count_1_io_out ? io_r_65_b : _GEN_644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_646 = 9'h42 == r_count_1_io_out ? io_r_66_b : _GEN_645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_647 = 9'h43 == r_count_1_io_out ? io_r_67_b : _GEN_646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_648 = 9'h44 == r_count_1_io_out ? io_r_68_b : _GEN_647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_649 = 9'h45 == r_count_1_io_out ? io_r_69_b : _GEN_648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_650 = 9'h46 == r_count_1_io_out ? io_r_70_b : _GEN_649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_651 = 9'h47 == r_count_1_io_out ? io_r_71_b : _GEN_650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_652 = 9'h48 == r_count_1_io_out ? io_r_72_b : _GEN_651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_653 = 9'h49 == r_count_1_io_out ? io_r_73_b : _GEN_652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_654 = 9'h4a == r_count_1_io_out ? io_r_74_b : _GEN_653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_655 = 9'h4b == r_count_1_io_out ? io_r_75_b : _GEN_654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_656 = 9'h4c == r_count_1_io_out ? io_r_76_b : _GEN_655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_657 = 9'h4d == r_count_1_io_out ? io_r_77_b : _GEN_656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_658 = 9'h4e == r_count_1_io_out ? io_r_78_b : _GEN_657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_659 = 9'h4f == r_count_1_io_out ? io_r_79_b : _GEN_658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_660 = 9'h50 == r_count_1_io_out ? io_r_80_b : _GEN_659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_661 = 9'h51 == r_count_1_io_out ? io_r_81_b : _GEN_660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_662 = 9'h52 == r_count_1_io_out ? io_r_82_b : _GEN_661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_663 = 9'h53 == r_count_1_io_out ? io_r_83_b : _GEN_662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_664 = 9'h54 == r_count_1_io_out ? io_r_84_b : _GEN_663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_665 = 9'h55 == r_count_1_io_out ? io_r_85_b : _GEN_664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_666 = 9'h56 == r_count_1_io_out ? io_r_86_b : _GEN_665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_667 = 9'h57 == r_count_1_io_out ? io_r_87_b : _GEN_666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_668 = 9'h58 == r_count_1_io_out ? io_r_88_b : _GEN_667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_669 = 9'h59 == r_count_1_io_out ? io_r_89_b : _GEN_668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_670 = 9'h5a == r_count_1_io_out ? io_r_90_b : _GEN_669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_671 = 9'h5b == r_count_1_io_out ? io_r_91_b : _GEN_670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_672 = 9'h5c == r_count_1_io_out ? io_r_92_b : _GEN_671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_673 = 9'h5d == r_count_1_io_out ? io_r_93_b : _GEN_672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_674 = 9'h5e == r_count_1_io_out ? io_r_94_b : _GEN_673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_675 = 9'h5f == r_count_1_io_out ? io_r_95_b : _GEN_674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_676 = 9'h60 == r_count_1_io_out ? io_r_96_b : _GEN_675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_677 = 9'h61 == r_count_1_io_out ? io_r_97_b : _GEN_676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_678 = 9'h62 == r_count_1_io_out ? io_r_98_b : _GEN_677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_679 = 9'h63 == r_count_1_io_out ? io_r_99_b : _GEN_678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_680 = 9'h64 == r_count_1_io_out ? io_r_100_b : _GEN_679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_681 = 9'h65 == r_count_1_io_out ? io_r_101_b : _GEN_680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_682 = 9'h66 == r_count_1_io_out ? io_r_102_b : _GEN_681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_683 = 9'h67 == r_count_1_io_out ? io_r_103_b : _GEN_682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_684 = 9'h68 == r_count_1_io_out ? io_r_104_b : _GEN_683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_685 = 9'h69 == r_count_1_io_out ? io_r_105_b : _GEN_684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_686 = 9'h6a == r_count_1_io_out ? io_r_106_b : _GEN_685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_687 = 9'h6b == r_count_1_io_out ? io_r_107_b : _GEN_686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_688 = 9'h6c == r_count_1_io_out ? io_r_108_b : _GEN_687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_689 = 9'h6d == r_count_1_io_out ? io_r_109_b : _GEN_688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_690 = 9'h6e == r_count_1_io_out ? io_r_110_b : _GEN_689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_691 = 9'h6f == r_count_1_io_out ? io_r_111_b : _GEN_690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_692 = 9'h70 == r_count_1_io_out ? io_r_112_b : _GEN_691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_693 = 9'h71 == r_count_1_io_out ? io_r_113_b : _GEN_692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_694 = 9'h72 == r_count_1_io_out ? io_r_114_b : _GEN_693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_695 = 9'h73 == r_count_1_io_out ? io_r_115_b : _GEN_694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_696 = 9'h74 == r_count_1_io_out ? io_r_116_b : _GEN_695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_697 = 9'h75 == r_count_1_io_out ? io_r_117_b : _GEN_696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_698 = 9'h76 == r_count_1_io_out ? io_r_118_b : _GEN_697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_699 = 9'h77 == r_count_1_io_out ? io_r_119_b : _GEN_698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_700 = 9'h78 == r_count_1_io_out ? io_r_120_b : _GEN_699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_701 = 9'h79 == r_count_1_io_out ? io_r_121_b : _GEN_700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_702 = 9'h7a == r_count_1_io_out ? io_r_122_b : _GEN_701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_703 = 9'h7b == r_count_1_io_out ? io_r_123_b : _GEN_702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_704 = 9'h7c == r_count_1_io_out ? io_r_124_b : _GEN_703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_705 = 9'h7d == r_count_1_io_out ? io_r_125_b : _GEN_704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_706 = 9'h7e == r_count_1_io_out ? io_r_126_b : _GEN_705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_707 = 9'h7f == r_count_1_io_out ? io_r_127_b : _GEN_706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_708 = 9'h80 == r_count_1_io_out ? io_r_128_b : _GEN_707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_709 = 9'h81 == r_count_1_io_out ? io_r_129_b : _GEN_708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_710 = 9'h82 == r_count_1_io_out ? io_r_130_b : _GEN_709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_711 = 9'h83 == r_count_1_io_out ? io_r_131_b : _GEN_710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_712 = 9'h84 == r_count_1_io_out ? io_r_132_b : _GEN_711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_713 = 9'h85 == r_count_1_io_out ? io_r_133_b : _GEN_712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_714 = 9'h86 == r_count_1_io_out ? io_r_134_b : _GEN_713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_715 = 9'h87 == r_count_1_io_out ? io_r_135_b : _GEN_714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_716 = 9'h88 == r_count_1_io_out ? io_r_136_b : _GEN_715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_717 = 9'h89 == r_count_1_io_out ? io_r_137_b : _GEN_716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_718 = 9'h8a == r_count_1_io_out ? io_r_138_b : _GEN_717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_719 = 9'h8b == r_count_1_io_out ? io_r_139_b : _GEN_718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_720 = 9'h8c == r_count_1_io_out ? io_r_140_b : _GEN_719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_721 = 9'h8d == r_count_1_io_out ? io_r_141_b : _GEN_720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_722 = 9'h8e == r_count_1_io_out ? io_r_142_b : _GEN_721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_723 = 9'h8f == r_count_1_io_out ? io_r_143_b : _GEN_722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_724 = 9'h90 == r_count_1_io_out ? io_r_144_b : _GEN_723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_725 = 9'h91 == r_count_1_io_out ? io_r_145_b : _GEN_724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_726 = 9'h92 == r_count_1_io_out ? io_r_146_b : _GEN_725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_727 = 9'h93 == r_count_1_io_out ? io_r_147_b : _GEN_726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_728 = 9'h94 == r_count_1_io_out ? io_r_148_b : _GEN_727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_729 = 9'h95 == r_count_1_io_out ? io_r_149_b : _GEN_728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_730 = 9'h96 == r_count_1_io_out ? io_r_150_b : _GEN_729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_731 = 9'h97 == r_count_1_io_out ? io_r_151_b : _GEN_730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_732 = 9'h98 == r_count_1_io_out ? io_r_152_b : _GEN_731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_733 = 9'h99 == r_count_1_io_out ? io_r_153_b : _GEN_732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_734 = 9'h9a == r_count_1_io_out ? io_r_154_b : _GEN_733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_735 = 9'h9b == r_count_1_io_out ? io_r_155_b : _GEN_734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_736 = 9'h9c == r_count_1_io_out ? io_r_156_b : _GEN_735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_737 = 9'h9d == r_count_1_io_out ? io_r_157_b : _GEN_736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_738 = 9'h9e == r_count_1_io_out ? io_r_158_b : _GEN_737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_739 = 9'h9f == r_count_1_io_out ? io_r_159_b : _GEN_738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_740 = 9'ha0 == r_count_1_io_out ? io_r_160_b : _GEN_739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_741 = 9'ha1 == r_count_1_io_out ? io_r_161_b : _GEN_740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_742 = 9'ha2 == r_count_1_io_out ? io_r_162_b : _GEN_741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_743 = 9'ha3 == r_count_1_io_out ? io_r_163_b : _GEN_742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_744 = 9'ha4 == r_count_1_io_out ? io_r_164_b : _GEN_743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_745 = 9'ha5 == r_count_1_io_out ? io_r_165_b : _GEN_744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_746 = 9'ha6 == r_count_1_io_out ? io_r_166_b : _GEN_745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_747 = 9'ha7 == r_count_1_io_out ? io_r_167_b : _GEN_746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_748 = 9'ha8 == r_count_1_io_out ? io_r_168_b : _GEN_747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_749 = 9'ha9 == r_count_1_io_out ? io_r_169_b : _GEN_748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_750 = 9'haa == r_count_1_io_out ? io_r_170_b : _GEN_749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_751 = 9'hab == r_count_1_io_out ? io_r_171_b : _GEN_750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_752 = 9'hac == r_count_1_io_out ? io_r_172_b : _GEN_751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_753 = 9'had == r_count_1_io_out ? io_r_173_b : _GEN_752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_754 = 9'hae == r_count_1_io_out ? io_r_174_b : _GEN_753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_755 = 9'haf == r_count_1_io_out ? io_r_175_b : _GEN_754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_756 = 9'hb0 == r_count_1_io_out ? io_r_176_b : _GEN_755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_757 = 9'hb1 == r_count_1_io_out ? io_r_177_b : _GEN_756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_758 = 9'hb2 == r_count_1_io_out ? io_r_178_b : _GEN_757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_759 = 9'hb3 == r_count_1_io_out ? io_r_179_b : _GEN_758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_760 = 9'hb4 == r_count_1_io_out ? io_r_180_b : _GEN_759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_761 = 9'hb5 == r_count_1_io_out ? io_r_181_b : _GEN_760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_762 = 9'hb6 == r_count_1_io_out ? io_r_182_b : _GEN_761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_763 = 9'hb7 == r_count_1_io_out ? io_r_183_b : _GEN_762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_764 = 9'hb8 == r_count_1_io_out ? io_r_184_b : _GEN_763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_765 = 9'hb9 == r_count_1_io_out ? io_r_185_b : _GEN_764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_766 = 9'hba == r_count_1_io_out ? io_r_186_b : _GEN_765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_767 = 9'hbb == r_count_1_io_out ? io_r_187_b : _GEN_766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_768 = 9'hbc == r_count_1_io_out ? io_r_188_b : _GEN_767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_769 = 9'hbd == r_count_1_io_out ? io_r_189_b : _GEN_768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_770 = 9'hbe == r_count_1_io_out ? io_r_190_b : _GEN_769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_771 = 9'hbf == r_count_1_io_out ? io_r_191_b : _GEN_770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_772 = 9'hc0 == r_count_1_io_out ? io_r_192_b : _GEN_771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_773 = 9'hc1 == r_count_1_io_out ? io_r_193_b : _GEN_772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_774 = 9'hc2 == r_count_1_io_out ? io_r_194_b : _GEN_773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_775 = 9'hc3 == r_count_1_io_out ? io_r_195_b : _GEN_774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_776 = 9'hc4 == r_count_1_io_out ? io_r_196_b : _GEN_775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_777 = 9'hc5 == r_count_1_io_out ? io_r_197_b : _GEN_776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_778 = 9'hc6 == r_count_1_io_out ? io_r_198_b : _GEN_777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_779 = 9'hc7 == r_count_1_io_out ? io_r_199_b : _GEN_778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_780 = 9'hc8 == r_count_1_io_out ? io_r_200_b : _GEN_779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_781 = 9'hc9 == r_count_1_io_out ? io_r_201_b : _GEN_780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_782 = 9'hca == r_count_1_io_out ? io_r_202_b : _GEN_781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_783 = 9'hcb == r_count_1_io_out ? io_r_203_b : _GEN_782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_784 = 9'hcc == r_count_1_io_out ? io_r_204_b : _GEN_783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_785 = 9'hcd == r_count_1_io_out ? io_r_205_b : _GEN_784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_786 = 9'hce == r_count_1_io_out ? io_r_206_b : _GEN_785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_787 = 9'hcf == r_count_1_io_out ? io_r_207_b : _GEN_786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_788 = 9'hd0 == r_count_1_io_out ? io_r_208_b : _GEN_787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_789 = 9'hd1 == r_count_1_io_out ? io_r_209_b : _GEN_788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_790 = 9'hd2 == r_count_1_io_out ? io_r_210_b : _GEN_789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_791 = 9'hd3 == r_count_1_io_out ? io_r_211_b : _GEN_790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_792 = 9'hd4 == r_count_1_io_out ? io_r_212_b : _GEN_791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_793 = 9'hd5 == r_count_1_io_out ? io_r_213_b : _GEN_792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_794 = 9'hd6 == r_count_1_io_out ? io_r_214_b : _GEN_793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_795 = 9'hd7 == r_count_1_io_out ? io_r_215_b : _GEN_794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_796 = 9'hd8 == r_count_1_io_out ? io_r_216_b : _GEN_795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_797 = 9'hd9 == r_count_1_io_out ? io_r_217_b : _GEN_796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_798 = 9'hda == r_count_1_io_out ? io_r_218_b : _GEN_797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_799 = 9'hdb == r_count_1_io_out ? io_r_219_b : _GEN_798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_800 = 9'hdc == r_count_1_io_out ? io_r_220_b : _GEN_799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_801 = 9'hdd == r_count_1_io_out ? io_r_221_b : _GEN_800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_802 = 9'hde == r_count_1_io_out ? io_r_222_b : _GEN_801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_803 = 9'hdf == r_count_1_io_out ? io_r_223_b : _GEN_802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_804 = 9'he0 == r_count_1_io_out ? io_r_224_b : _GEN_803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_805 = 9'he1 == r_count_1_io_out ? io_r_225_b : _GEN_804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_806 = 9'he2 == r_count_1_io_out ? io_r_226_b : _GEN_805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_807 = 9'he3 == r_count_1_io_out ? io_r_227_b : _GEN_806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_808 = 9'he4 == r_count_1_io_out ? io_r_228_b : _GEN_807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_809 = 9'he5 == r_count_1_io_out ? io_r_229_b : _GEN_808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_810 = 9'he6 == r_count_1_io_out ? io_r_230_b : _GEN_809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_811 = 9'he7 == r_count_1_io_out ? io_r_231_b : _GEN_810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_812 = 9'he8 == r_count_1_io_out ? io_r_232_b : _GEN_811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_813 = 9'he9 == r_count_1_io_out ? io_r_233_b : _GEN_812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_814 = 9'hea == r_count_1_io_out ? io_r_234_b : _GEN_813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_815 = 9'heb == r_count_1_io_out ? io_r_235_b : _GEN_814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_816 = 9'hec == r_count_1_io_out ? io_r_236_b : _GEN_815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_817 = 9'hed == r_count_1_io_out ? io_r_237_b : _GEN_816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_818 = 9'hee == r_count_1_io_out ? io_r_238_b : _GEN_817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_819 = 9'hef == r_count_1_io_out ? io_r_239_b : _GEN_818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_820 = 9'hf0 == r_count_1_io_out ? io_r_240_b : _GEN_819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_821 = 9'hf1 == r_count_1_io_out ? io_r_241_b : _GEN_820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_822 = 9'hf2 == r_count_1_io_out ? io_r_242_b : _GEN_821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_823 = 9'hf3 == r_count_1_io_out ? io_r_243_b : _GEN_822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_824 = 9'hf4 == r_count_1_io_out ? io_r_244_b : _GEN_823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_825 = 9'hf5 == r_count_1_io_out ? io_r_245_b : _GEN_824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_826 = 9'hf6 == r_count_1_io_out ? io_r_246_b : _GEN_825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_827 = 9'hf7 == r_count_1_io_out ? io_r_247_b : _GEN_826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_828 = 9'hf8 == r_count_1_io_out ? io_r_248_b : _GEN_827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_829 = 9'hf9 == r_count_1_io_out ? io_r_249_b : _GEN_828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_830 = 9'hfa == r_count_1_io_out ? io_r_250_b : _GEN_829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_831 = 9'hfb == r_count_1_io_out ? io_r_251_b : _GEN_830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_832 = 9'hfc == r_count_1_io_out ? io_r_252_b : _GEN_831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_833 = 9'hfd == r_count_1_io_out ? io_r_253_b : _GEN_832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_834 = 9'hfe == r_count_1_io_out ? io_r_254_b : _GEN_833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_835 = 9'hff == r_count_1_io_out ? io_r_255_b : _GEN_834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_836 = 9'h100 == r_count_1_io_out ? io_r_256_b : _GEN_835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_837 = 9'h101 == r_count_1_io_out ? io_r_257_b : _GEN_836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_838 = 9'h102 == r_count_1_io_out ? io_r_258_b : _GEN_837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_839 = 9'h103 == r_count_1_io_out ? io_r_259_b : _GEN_838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_840 = 9'h104 == r_count_1_io_out ? io_r_260_b : _GEN_839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_841 = 9'h105 == r_count_1_io_out ? io_r_261_b : _GEN_840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_842 = 9'h106 == r_count_1_io_out ? io_r_262_b : _GEN_841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_843 = 9'h107 == r_count_1_io_out ? io_r_263_b : _GEN_842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_844 = 9'h108 == r_count_1_io_out ? io_r_264_b : _GEN_843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_845 = 9'h109 == r_count_1_io_out ? io_r_265_b : _GEN_844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_846 = 9'h10a == r_count_1_io_out ? io_r_266_b : _GEN_845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_847 = 9'h10b == r_count_1_io_out ? io_r_267_b : _GEN_846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_848 = 9'h10c == r_count_1_io_out ? io_r_268_b : _GEN_847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_849 = 9'h10d == r_count_1_io_out ? io_r_269_b : _GEN_848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_850 = 9'h10e == r_count_1_io_out ? io_r_270_b : _GEN_849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_851 = 9'h10f == r_count_1_io_out ? io_r_271_b : _GEN_850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_852 = 9'h110 == r_count_1_io_out ? io_r_272_b : _GEN_851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_853 = 9'h111 == r_count_1_io_out ? io_r_273_b : _GEN_852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_854 = 9'h112 == r_count_1_io_out ? io_r_274_b : _GEN_853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_855 = 9'h113 == r_count_1_io_out ? io_r_275_b : _GEN_854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_856 = 9'h114 == r_count_1_io_out ? io_r_276_b : _GEN_855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_857 = 9'h115 == r_count_1_io_out ? io_r_277_b : _GEN_856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_858 = 9'h116 == r_count_1_io_out ? io_r_278_b : _GEN_857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_859 = 9'h117 == r_count_1_io_out ? io_r_279_b : _GEN_858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_860 = 9'h118 == r_count_1_io_out ? io_r_280_b : _GEN_859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_861 = 9'h119 == r_count_1_io_out ? io_r_281_b : _GEN_860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_862 = 9'h11a == r_count_1_io_out ? io_r_282_b : _GEN_861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_863 = 9'h11b == r_count_1_io_out ? io_r_283_b : _GEN_862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_864 = 9'h11c == r_count_1_io_out ? io_r_284_b : _GEN_863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_865 = 9'h11d == r_count_1_io_out ? io_r_285_b : _GEN_864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_866 = 9'h11e == r_count_1_io_out ? io_r_286_b : _GEN_865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_867 = 9'h11f == r_count_1_io_out ? io_r_287_b : _GEN_866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_868 = 9'h120 == r_count_1_io_out ? io_r_288_b : _GEN_867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_869 = 9'h121 == r_count_1_io_out ? io_r_289_b : _GEN_868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_870 = 9'h122 == r_count_1_io_out ? io_r_290_b : _GEN_869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_871 = 9'h123 == r_count_1_io_out ? io_r_291_b : _GEN_870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_872 = 9'h124 == r_count_1_io_out ? io_r_292_b : _GEN_871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_873 = 9'h125 == r_count_1_io_out ? io_r_293_b : _GEN_872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_874 = 9'h126 == r_count_1_io_out ? io_r_294_b : _GEN_873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_875 = 9'h127 == r_count_1_io_out ? io_r_295_b : _GEN_874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_876 = 9'h128 == r_count_1_io_out ? io_r_296_b : _GEN_875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_877 = 9'h129 == r_count_1_io_out ? io_r_297_b : _GEN_876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_878 = 9'h12a == r_count_1_io_out ? io_r_298_b : _GEN_877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_879 = 9'h12b == r_count_1_io_out ? io_r_299_b : _GEN_878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_880 = 9'h12c == r_count_1_io_out ? io_r_300_b : _GEN_879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_881 = 9'h12d == r_count_1_io_out ? io_r_301_b : _GEN_880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_882 = 9'h12e == r_count_1_io_out ? io_r_302_b : _GEN_881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_883 = 9'h12f == r_count_1_io_out ? io_r_303_b : _GEN_882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_884 = 9'h130 == r_count_1_io_out ? io_r_304_b : _GEN_883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_885 = 9'h131 == r_count_1_io_out ? io_r_305_b : _GEN_884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_886 = 9'h132 == r_count_1_io_out ? io_r_306_b : _GEN_885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_887 = 9'h133 == r_count_1_io_out ? io_r_307_b : _GEN_886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_888 = 9'h134 == r_count_1_io_out ? io_r_308_b : _GEN_887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_889 = 9'h135 == r_count_1_io_out ? io_r_309_b : _GEN_888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_890 = 9'h136 == r_count_1_io_out ? io_r_310_b : _GEN_889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_891 = 9'h137 == r_count_1_io_out ? io_r_311_b : _GEN_890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_892 = 9'h138 == r_count_1_io_out ? io_r_312_b : _GEN_891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_893 = 9'h139 == r_count_1_io_out ? io_r_313_b : _GEN_892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_894 = 9'h13a == r_count_1_io_out ? io_r_314_b : _GEN_893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_895 = 9'h13b == r_count_1_io_out ? io_r_315_b : _GEN_894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_896 = 9'h13c == r_count_1_io_out ? io_r_316_b : _GEN_895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_897 = 9'h13d == r_count_1_io_out ? io_r_317_b : _GEN_896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_898 = 9'h13e == r_count_1_io_out ? io_r_318_b : _GEN_897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_899 = 9'h13f == r_count_1_io_out ? io_r_319_b : _GEN_898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_900 = 9'h140 == r_count_1_io_out ? io_r_320_b : _GEN_899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_901 = 9'h141 == r_count_1_io_out ? io_r_321_b : _GEN_900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_902 = 9'h142 == r_count_1_io_out ? io_r_322_b : _GEN_901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_903 = 9'h143 == r_count_1_io_out ? io_r_323_b : _GEN_902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_904 = 9'h144 == r_count_1_io_out ? io_r_324_b : _GEN_903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_905 = 9'h145 == r_count_1_io_out ? io_r_325_b : _GEN_904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_906 = 9'h146 == r_count_1_io_out ? io_r_326_b : _GEN_905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_907 = 9'h147 == r_count_1_io_out ? io_r_327_b : _GEN_906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_908 = 9'h148 == r_count_1_io_out ? io_r_328_b : _GEN_907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_909 = 9'h149 == r_count_1_io_out ? io_r_329_b : _GEN_908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_910 = 9'h14a == r_count_1_io_out ? io_r_330_b : _GEN_909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_911 = 9'h14b == r_count_1_io_out ? io_r_331_b : _GEN_910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_912 = 9'h14c == r_count_1_io_out ? io_r_332_b : _GEN_911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_913 = 9'h14d == r_count_1_io_out ? io_r_333_b : _GEN_912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_914 = 9'h14e == r_count_1_io_out ? io_r_334_b : _GEN_913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_915 = 9'h14f == r_count_1_io_out ? io_r_335_b : _GEN_914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_916 = 9'h150 == r_count_1_io_out ? io_r_336_b : _GEN_915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_917 = 9'h151 == r_count_1_io_out ? io_r_337_b : _GEN_916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_918 = 9'h152 == r_count_1_io_out ? io_r_338_b : _GEN_917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_919 = 9'h153 == r_count_1_io_out ? io_r_339_b : _GEN_918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_920 = 9'h154 == r_count_1_io_out ? io_r_340_b : _GEN_919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_921 = 9'h155 == r_count_1_io_out ? io_r_341_b : _GEN_920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_922 = 9'h156 == r_count_1_io_out ? io_r_342_b : _GEN_921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_923 = 9'h157 == r_count_1_io_out ? io_r_343_b : _GEN_922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_924 = 9'h158 == r_count_1_io_out ? io_r_344_b : _GEN_923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_925 = 9'h159 == r_count_1_io_out ? io_r_345_b : _GEN_924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_926 = 9'h15a == r_count_1_io_out ? io_r_346_b : _GEN_925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_927 = 9'h15b == r_count_1_io_out ? io_r_347_b : _GEN_926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_928 = 9'h15c == r_count_1_io_out ? io_r_348_b : _GEN_927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_929 = 9'h15d == r_count_1_io_out ? io_r_349_b : _GEN_928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_930 = 9'h15e == r_count_1_io_out ? io_r_350_b : _GEN_929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_931 = 9'h15f == r_count_1_io_out ? io_r_351_b : _GEN_930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_932 = 9'h160 == r_count_1_io_out ? io_r_352_b : _GEN_931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_933 = 9'h161 == r_count_1_io_out ? io_r_353_b : _GEN_932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_934 = 9'h162 == r_count_1_io_out ? io_r_354_b : _GEN_933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_935 = 9'h163 == r_count_1_io_out ? io_r_355_b : _GEN_934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_936 = 9'h164 == r_count_1_io_out ? io_r_356_b : _GEN_935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_937 = 9'h165 == r_count_1_io_out ? io_r_357_b : _GEN_936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_938 = 9'h166 == r_count_1_io_out ? io_r_358_b : _GEN_937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_939 = 9'h167 == r_count_1_io_out ? io_r_359_b : _GEN_938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_940 = 9'h168 == r_count_1_io_out ? io_r_360_b : _GEN_939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_941 = 9'h169 == r_count_1_io_out ? io_r_361_b : _GEN_940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_942 = 9'h16a == r_count_1_io_out ? io_r_362_b : _GEN_941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_943 = 9'h16b == r_count_1_io_out ? io_r_363_b : _GEN_942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_944 = 9'h16c == r_count_1_io_out ? io_r_364_b : _GEN_943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_945 = 9'h16d == r_count_1_io_out ? io_r_365_b : _GEN_944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_946 = 9'h16e == r_count_1_io_out ? io_r_366_b : _GEN_945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_947 = 9'h16f == r_count_1_io_out ? io_r_367_b : _GEN_946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_948 = 9'h170 == r_count_1_io_out ? io_r_368_b : _GEN_947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_949 = 9'h171 == r_count_1_io_out ? io_r_369_b : _GEN_948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_950 = 9'h172 == r_count_1_io_out ? io_r_370_b : _GEN_949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_951 = 9'h173 == r_count_1_io_out ? io_r_371_b : _GEN_950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_952 = 9'h174 == r_count_1_io_out ? io_r_372_b : _GEN_951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_953 = 9'h175 == r_count_1_io_out ? io_r_373_b : _GEN_952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_954 = 9'h176 == r_count_1_io_out ? io_r_374_b : _GEN_953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_955 = 9'h177 == r_count_1_io_out ? io_r_375_b : _GEN_954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_956 = 9'h178 == r_count_1_io_out ? io_r_376_b : _GEN_955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_957 = 9'h179 == r_count_1_io_out ? io_r_377_b : _GEN_956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_958 = 9'h17a == r_count_1_io_out ? io_r_378_b : _GEN_957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_959 = 9'h17b == r_count_1_io_out ? io_r_379_b : _GEN_958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_960 = 9'h17c == r_count_1_io_out ? io_r_380_b : _GEN_959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_961 = 9'h17d == r_count_1_io_out ? io_r_381_b : _GEN_960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_962 = 9'h17e == r_count_1_io_out ? io_r_382_b : _GEN_961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_963 = 9'h17f == r_count_1_io_out ? io_r_383_b : _GEN_962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_964 = 9'h180 == r_count_1_io_out ? io_r_384_b : _GEN_963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_965 = 9'h181 == r_count_1_io_out ? io_r_385_b : _GEN_964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_966 = 9'h182 == r_count_1_io_out ? io_r_386_b : _GEN_965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_967 = 9'h183 == r_count_1_io_out ? io_r_387_b : _GEN_966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_968 = 9'h184 == r_count_1_io_out ? io_r_388_b : _GEN_967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_969 = 9'h185 == r_count_1_io_out ? io_r_389_b : _GEN_968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_970 = 9'h186 == r_count_1_io_out ? io_r_390_b : _GEN_969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_971 = 9'h187 == r_count_1_io_out ? io_r_391_b : _GEN_970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_972 = 9'h188 == r_count_1_io_out ? io_r_392_b : _GEN_971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_973 = 9'h189 == r_count_1_io_out ? io_r_393_b : _GEN_972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_974 = 9'h18a == r_count_1_io_out ? io_r_394_b : _GEN_973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_975 = 9'h18b == r_count_1_io_out ? io_r_395_b : _GEN_974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_976 = 9'h18c == r_count_1_io_out ? io_r_396_b : _GEN_975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_977 = 9'h18d == r_count_1_io_out ? io_r_397_b : _GEN_976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_978 = 9'h18e == r_count_1_io_out ? io_r_398_b : _GEN_977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_981 = 9'h1 == r_count_2_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_982 = 9'h2 == r_count_2_io_out ? io_r_2_b : _GEN_981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_983 = 9'h3 == r_count_2_io_out ? io_r_3_b : _GEN_982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_984 = 9'h4 == r_count_2_io_out ? io_r_4_b : _GEN_983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_985 = 9'h5 == r_count_2_io_out ? io_r_5_b : _GEN_984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_986 = 9'h6 == r_count_2_io_out ? io_r_6_b : _GEN_985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_987 = 9'h7 == r_count_2_io_out ? io_r_7_b : _GEN_986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_988 = 9'h8 == r_count_2_io_out ? io_r_8_b : _GEN_987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_989 = 9'h9 == r_count_2_io_out ? io_r_9_b : _GEN_988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_990 = 9'ha == r_count_2_io_out ? io_r_10_b : _GEN_989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_991 = 9'hb == r_count_2_io_out ? io_r_11_b : _GEN_990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_992 = 9'hc == r_count_2_io_out ? io_r_12_b : _GEN_991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_993 = 9'hd == r_count_2_io_out ? io_r_13_b : _GEN_992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_994 = 9'he == r_count_2_io_out ? io_r_14_b : _GEN_993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_995 = 9'hf == r_count_2_io_out ? io_r_15_b : _GEN_994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_996 = 9'h10 == r_count_2_io_out ? io_r_16_b : _GEN_995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_997 = 9'h11 == r_count_2_io_out ? io_r_17_b : _GEN_996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_998 = 9'h12 == r_count_2_io_out ? io_r_18_b : _GEN_997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_999 = 9'h13 == r_count_2_io_out ? io_r_19_b : _GEN_998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1000 = 9'h14 == r_count_2_io_out ? io_r_20_b : _GEN_999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1001 = 9'h15 == r_count_2_io_out ? io_r_21_b : _GEN_1000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1002 = 9'h16 == r_count_2_io_out ? io_r_22_b : _GEN_1001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1003 = 9'h17 == r_count_2_io_out ? io_r_23_b : _GEN_1002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1004 = 9'h18 == r_count_2_io_out ? io_r_24_b : _GEN_1003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1005 = 9'h19 == r_count_2_io_out ? io_r_25_b : _GEN_1004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1006 = 9'h1a == r_count_2_io_out ? io_r_26_b : _GEN_1005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1007 = 9'h1b == r_count_2_io_out ? io_r_27_b : _GEN_1006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1008 = 9'h1c == r_count_2_io_out ? io_r_28_b : _GEN_1007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1009 = 9'h1d == r_count_2_io_out ? io_r_29_b : _GEN_1008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1010 = 9'h1e == r_count_2_io_out ? io_r_30_b : _GEN_1009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1011 = 9'h1f == r_count_2_io_out ? io_r_31_b : _GEN_1010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1012 = 9'h20 == r_count_2_io_out ? io_r_32_b : _GEN_1011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1013 = 9'h21 == r_count_2_io_out ? io_r_33_b : _GEN_1012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1014 = 9'h22 == r_count_2_io_out ? io_r_34_b : _GEN_1013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1015 = 9'h23 == r_count_2_io_out ? io_r_35_b : _GEN_1014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1016 = 9'h24 == r_count_2_io_out ? io_r_36_b : _GEN_1015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1017 = 9'h25 == r_count_2_io_out ? io_r_37_b : _GEN_1016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1018 = 9'h26 == r_count_2_io_out ? io_r_38_b : _GEN_1017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1019 = 9'h27 == r_count_2_io_out ? io_r_39_b : _GEN_1018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1020 = 9'h28 == r_count_2_io_out ? io_r_40_b : _GEN_1019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1021 = 9'h29 == r_count_2_io_out ? io_r_41_b : _GEN_1020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1022 = 9'h2a == r_count_2_io_out ? io_r_42_b : _GEN_1021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1023 = 9'h2b == r_count_2_io_out ? io_r_43_b : _GEN_1022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1024 = 9'h2c == r_count_2_io_out ? io_r_44_b : _GEN_1023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1025 = 9'h2d == r_count_2_io_out ? io_r_45_b : _GEN_1024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1026 = 9'h2e == r_count_2_io_out ? io_r_46_b : _GEN_1025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1027 = 9'h2f == r_count_2_io_out ? io_r_47_b : _GEN_1026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1028 = 9'h30 == r_count_2_io_out ? io_r_48_b : _GEN_1027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1029 = 9'h31 == r_count_2_io_out ? io_r_49_b : _GEN_1028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1030 = 9'h32 == r_count_2_io_out ? io_r_50_b : _GEN_1029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1031 = 9'h33 == r_count_2_io_out ? io_r_51_b : _GEN_1030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1032 = 9'h34 == r_count_2_io_out ? io_r_52_b : _GEN_1031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1033 = 9'h35 == r_count_2_io_out ? io_r_53_b : _GEN_1032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1034 = 9'h36 == r_count_2_io_out ? io_r_54_b : _GEN_1033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1035 = 9'h37 == r_count_2_io_out ? io_r_55_b : _GEN_1034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1036 = 9'h38 == r_count_2_io_out ? io_r_56_b : _GEN_1035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1037 = 9'h39 == r_count_2_io_out ? io_r_57_b : _GEN_1036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1038 = 9'h3a == r_count_2_io_out ? io_r_58_b : _GEN_1037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1039 = 9'h3b == r_count_2_io_out ? io_r_59_b : _GEN_1038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1040 = 9'h3c == r_count_2_io_out ? io_r_60_b : _GEN_1039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1041 = 9'h3d == r_count_2_io_out ? io_r_61_b : _GEN_1040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1042 = 9'h3e == r_count_2_io_out ? io_r_62_b : _GEN_1041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1043 = 9'h3f == r_count_2_io_out ? io_r_63_b : _GEN_1042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1044 = 9'h40 == r_count_2_io_out ? io_r_64_b : _GEN_1043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1045 = 9'h41 == r_count_2_io_out ? io_r_65_b : _GEN_1044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1046 = 9'h42 == r_count_2_io_out ? io_r_66_b : _GEN_1045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1047 = 9'h43 == r_count_2_io_out ? io_r_67_b : _GEN_1046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1048 = 9'h44 == r_count_2_io_out ? io_r_68_b : _GEN_1047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1049 = 9'h45 == r_count_2_io_out ? io_r_69_b : _GEN_1048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1050 = 9'h46 == r_count_2_io_out ? io_r_70_b : _GEN_1049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1051 = 9'h47 == r_count_2_io_out ? io_r_71_b : _GEN_1050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1052 = 9'h48 == r_count_2_io_out ? io_r_72_b : _GEN_1051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1053 = 9'h49 == r_count_2_io_out ? io_r_73_b : _GEN_1052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1054 = 9'h4a == r_count_2_io_out ? io_r_74_b : _GEN_1053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1055 = 9'h4b == r_count_2_io_out ? io_r_75_b : _GEN_1054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1056 = 9'h4c == r_count_2_io_out ? io_r_76_b : _GEN_1055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1057 = 9'h4d == r_count_2_io_out ? io_r_77_b : _GEN_1056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1058 = 9'h4e == r_count_2_io_out ? io_r_78_b : _GEN_1057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1059 = 9'h4f == r_count_2_io_out ? io_r_79_b : _GEN_1058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1060 = 9'h50 == r_count_2_io_out ? io_r_80_b : _GEN_1059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1061 = 9'h51 == r_count_2_io_out ? io_r_81_b : _GEN_1060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1062 = 9'h52 == r_count_2_io_out ? io_r_82_b : _GEN_1061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1063 = 9'h53 == r_count_2_io_out ? io_r_83_b : _GEN_1062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1064 = 9'h54 == r_count_2_io_out ? io_r_84_b : _GEN_1063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1065 = 9'h55 == r_count_2_io_out ? io_r_85_b : _GEN_1064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1066 = 9'h56 == r_count_2_io_out ? io_r_86_b : _GEN_1065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1067 = 9'h57 == r_count_2_io_out ? io_r_87_b : _GEN_1066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1068 = 9'h58 == r_count_2_io_out ? io_r_88_b : _GEN_1067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1069 = 9'h59 == r_count_2_io_out ? io_r_89_b : _GEN_1068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1070 = 9'h5a == r_count_2_io_out ? io_r_90_b : _GEN_1069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1071 = 9'h5b == r_count_2_io_out ? io_r_91_b : _GEN_1070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1072 = 9'h5c == r_count_2_io_out ? io_r_92_b : _GEN_1071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1073 = 9'h5d == r_count_2_io_out ? io_r_93_b : _GEN_1072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1074 = 9'h5e == r_count_2_io_out ? io_r_94_b : _GEN_1073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1075 = 9'h5f == r_count_2_io_out ? io_r_95_b : _GEN_1074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1076 = 9'h60 == r_count_2_io_out ? io_r_96_b : _GEN_1075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1077 = 9'h61 == r_count_2_io_out ? io_r_97_b : _GEN_1076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1078 = 9'h62 == r_count_2_io_out ? io_r_98_b : _GEN_1077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1079 = 9'h63 == r_count_2_io_out ? io_r_99_b : _GEN_1078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1080 = 9'h64 == r_count_2_io_out ? io_r_100_b : _GEN_1079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1081 = 9'h65 == r_count_2_io_out ? io_r_101_b : _GEN_1080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1082 = 9'h66 == r_count_2_io_out ? io_r_102_b : _GEN_1081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1083 = 9'h67 == r_count_2_io_out ? io_r_103_b : _GEN_1082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1084 = 9'h68 == r_count_2_io_out ? io_r_104_b : _GEN_1083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1085 = 9'h69 == r_count_2_io_out ? io_r_105_b : _GEN_1084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1086 = 9'h6a == r_count_2_io_out ? io_r_106_b : _GEN_1085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1087 = 9'h6b == r_count_2_io_out ? io_r_107_b : _GEN_1086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1088 = 9'h6c == r_count_2_io_out ? io_r_108_b : _GEN_1087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1089 = 9'h6d == r_count_2_io_out ? io_r_109_b : _GEN_1088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1090 = 9'h6e == r_count_2_io_out ? io_r_110_b : _GEN_1089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1091 = 9'h6f == r_count_2_io_out ? io_r_111_b : _GEN_1090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1092 = 9'h70 == r_count_2_io_out ? io_r_112_b : _GEN_1091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1093 = 9'h71 == r_count_2_io_out ? io_r_113_b : _GEN_1092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1094 = 9'h72 == r_count_2_io_out ? io_r_114_b : _GEN_1093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1095 = 9'h73 == r_count_2_io_out ? io_r_115_b : _GEN_1094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1096 = 9'h74 == r_count_2_io_out ? io_r_116_b : _GEN_1095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1097 = 9'h75 == r_count_2_io_out ? io_r_117_b : _GEN_1096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1098 = 9'h76 == r_count_2_io_out ? io_r_118_b : _GEN_1097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1099 = 9'h77 == r_count_2_io_out ? io_r_119_b : _GEN_1098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1100 = 9'h78 == r_count_2_io_out ? io_r_120_b : _GEN_1099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1101 = 9'h79 == r_count_2_io_out ? io_r_121_b : _GEN_1100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1102 = 9'h7a == r_count_2_io_out ? io_r_122_b : _GEN_1101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1103 = 9'h7b == r_count_2_io_out ? io_r_123_b : _GEN_1102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1104 = 9'h7c == r_count_2_io_out ? io_r_124_b : _GEN_1103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1105 = 9'h7d == r_count_2_io_out ? io_r_125_b : _GEN_1104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1106 = 9'h7e == r_count_2_io_out ? io_r_126_b : _GEN_1105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1107 = 9'h7f == r_count_2_io_out ? io_r_127_b : _GEN_1106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1108 = 9'h80 == r_count_2_io_out ? io_r_128_b : _GEN_1107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1109 = 9'h81 == r_count_2_io_out ? io_r_129_b : _GEN_1108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1110 = 9'h82 == r_count_2_io_out ? io_r_130_b : _GEN_1109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1111 = 9'h83 == r_count_2_io_out ? io_r_131_b : _GEN_1110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1112 = 9'h84 == r_count_2_io_out ? io_r_132_b : _GEN_1111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1113 = 9'h85 == r_count_2_io_out ? io_r_133_b : _GEN_1112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1114 = 9'h86 == r_count_2_io_out ? io_r_134_b : _GEN_1113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1115 = 9'h87 == r_count_2_io_out ? io_r_135_b : _GEN_1114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1116 = 9'h88 == r_count_2_io_out ? io_r_136_b : _GEN_1115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1117 = 9'h89 == r_count_2_io_out ? io_r_137_b : _GEN_1116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1118 = 9'h8a == r_count_2_io_out ? io_r_138_b : _GEN_1117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1119 = 9'h8b == r_count_2_io_out ? io_r_139_b : _GEN_1118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1120 = 9'h8c == r_count_2_io_out ? io_r_140_b : _GEN_1119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1121 = 9'h8d == r_count_2_io_out ? io_r_141_b : _GEN_1120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1122 = 9'h8e == r_count_2_io_out ? io_r_142_b : _GEN_1121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1123 = 9'h8f == r_count_2_io_out ? io_r_143_b : _GEN_1122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1124 = 9'h90 == r_count_2_io_out ? io_r_144_b : _GEN_1123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1125 = 9'h91 == r_count_2_io_out ? io_r_145_b : _GEN_1124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1126 = 9'h92 == r_count_2_io_out ? io_r_146_b : _GEN_1125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1127 = 9'h93 == r_count_2_io_out ? io_r_147_b : _GEN_1126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1128 = 9'h94 == r_count_2_io_out ? io_r_148_b : _GEN_1127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1129 = 9'h95 == r_count_2_io_out ? io_r_149_b : _GEN_1128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1130 = 9'h96 == r_count_2_io_out ? io_r_150_b : _GEN_1129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1131 = 9'h97 == r_count_2_io_out ? io_r_151_b : _GEN_1130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1132 = 9'h98 == r_count_2_io_out ? io_r_152_b : _GEN_1131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1133 = 9'h99 == r_count_2_io_out ? io_r_153_b : _GEN_1132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1134 = 9'h9a == r_count_2_io_out ? io_r_154_b : _GEN_1133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1135 = 9'h9b == r_count_2_io_out ? io_r_155_b : _GEN_1134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1136 = 9'h9c == r_count_2_io_out ? io_r_156_b : _GEN_1135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1137 = 9'h9d == r_count_2_io_out ? io_r_157_b : _GEN_1136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1138 = 9'h9e == r_count_2_io_out ? io_r_158_b : _GEN_1137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1139 = 9'h9f == r_count_2_io_out ? io_r_159_b : _GEN_1138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1140 = 9'ha0 == r_count_2_io_out ? io_r_160_b : _GEN_1139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1141 = 9'ha1 == r_count_2_io_out ? io_r_161_b : _GEN_1140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1142 = 9'ha2 == r_count_2_io_out ? io_r_162_b : _GEN_1141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1143 = 9'ha3 == r_count_2_io_out ? io_r_163_b : _GEN_1142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1144 = 9'ha4 == r_count_2_io_out ? io_r_164_b : _GEN_1143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1145 = 9'ha5 == r_count_2_io_out ? io_r_165_b : _GEN_1144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1146 = 9'ha6 == r_count_2_io_out ? io_r_166_b : _GEN_1145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1147 = 9'ha7 == r_count_2_io_out ? io_r_167_b : _GEN_1146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1148 = 9'ha8 == r_count_2_io_out ? io_r_168_b : _GEN_1147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1149 = 9'ha9 == r_count_2_io_out ? io_r_169_b : _GEN_1148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1150 = 9'haa == r_count_2_io_out ? io_r_170_b : _GEN_1149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1151 = 9'hab == r_count_2_io_out ? io_r_171_b : _GEN_1150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1152 = 9'hac == r_count_2_io_out ? io_r_172_b : _GEN_1151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1153 = 9'had == r_count_2_io_out ? io_r_173_b : _GEN_1152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1154 = 9'hae == r_count_2_io_out ? io_r_174_b : _GEN_1153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1155 = 9'haf == r_count_2_io_out ? io_r_175_b : _GEN_1154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1156 = 9'hb0 == r_count_2_io_out ? io_r_176_b : _GEN_1155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1157 = 9'hb1 == r_count_2_io_out ? io_r_177_b : _GEN_1156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1158 = 9'hb2 == r_count_2_io_out ? io_r_178_b : _GEN_1157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1159 = 9'hb3 == r_count_2_io_out ? io_r_179_b : _GEN_1158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1160 = 9'hb4 == r_count_2_io_out ? io_r_180_b : _GEN_1159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1161 = 9'hb5 == r_count_2_io_out ? io_r_181_b : _GEN_1160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1162 = 9'hb6 == r_count_2_io_out ? io_r_182_b : _GEN_1161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1163 = 9'hb7 == r_count_2_io_out ? io_r_183_b : _GEN_1162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1164 = 9'hb8 == r_count_2_io_out ? io_r_184_b : _GEN_1163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1165 = 9'hb9 == r_count_2_io_out ? io_r_185_b : _GEN_1164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1166 = 9'hba == r_count_2_io_out ? io_r_186_b : _GEN_1165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1167 = 9'hbb == r_count_2_io_out ? io_r_187_b : _GEN_1166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1168 = 9'hbc == r_count_2_io_out ? io_r_188_b : _GEN_1167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1169 = 9'hbd == r_count_2_io_out ? io_r_189_b : _GEN_1168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1170 = 9'hbe == r_count_2_io_out ? io_r_190_b : _GEN_1169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1171 = 9'hbf == r_count_2_io_out ? io_r_191_b : _GEN_1170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1172 = 9'hc0 == r_count_2_io_out ? io_r_192_b : _GEN_1171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1173 = 9'hc1 == r_count_2_io_out ? io_r_193_b : _GEN_1172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1174 = 9'hc2 == r_count_2_io_out ? io_r_194_b : _GEN_1173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1175 = 9'hc3 == r_count_2_io_out ? io_r_195_b : _GEN_1174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1176 = 9'hc4 == r_count_2_io_out ? io_r_196_b : _GEN_1175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1177 = 9'hc5 == r_count_2_io_out ? io_r_197_b : _GEN_1176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1178 = 9'hc6 == r_count_2_io_out ? io_r_198_b : _GEN_1177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1179 = 9'hc7 == r_count_2_io_out ? io_r_199_b : _GEN_1178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1180 = 9'hc8 == r_count_2_io_out ? io_r_200_b : _GEN_1179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1181 = 9'hc9 == r_count_2_io_out ? io_r_201_b : _GEN_1180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1182 = 9'hca == r_count_2_io_out ? io_r_202_b : _GEN_1181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1183 = 9'hcb == r_count_2_io_out ? io_r_203_b : _GEN_1182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1184 = 9'hcc == r_count_2_io_out ? io_r_204_b : _GEN_1183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1185 = 9'hcd == r_count_2_io_out ? io_r_205_b : _GEN_1184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1186 = 9'hce == r_count_2_io_out ? io_r_206_b : _GEN_1185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1187 = 9'hcf == r_count_2_io_out ? io_r_207_b : _GEN_1186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1188 = 9'hd0 == r_count_2_io_out ? io_r_208_b : _GEN_1187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1189 = 9'hd1 == r_count_2_io_out ? io_r_209_b : _GEN_1188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1190 = 9'hd2 == r_count_2_io_out ? io_r_210_b : _GEN_1189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1191 = 9'hd3 == r_count_2_io_out ? io_r_211_b : _GEN_1190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1192 = 9'hd4 == r_count_2_io_out ? io_r_212_b : _GEN_1191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1193 = 9'hd5 == r_count_2_io_out ? io_r_213_b : _GEN_1192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1194 = 9'hd6 == r_count_2_io_out ? io_r_214_b : _GEN_1193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1195 = 9'hd7 == r_count_2_io_out ? io_r_215_b : _GEN_1194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1196 = 9'hd8 == r_count_2_io_out ? io_r_216_b : _GEN_1195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1197 = 9'hd9 == r_count_2_io_out ? io_r_217_b : _GEN_1196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1198 = 9'hda == r_count_2_io_out ? io_r_218_b : _GEN_1197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1199 = 9'hdb == r_count_2_io_out ? io_r_219_b : _GEN_1198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1200 = 9'hdc == r_count_2_io_out ? io_r_220_b : _GEN_1199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1201 = 9'hdd == r_count_2_io_out ? io_r_221_b : _GEN_1200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1202 = 9'hde == r_count_2_io_out ? io_r_222_b : _GEN_1201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1203 = 9'hdf == r_count_2_io_out ? io_r_223_b : _GEN_1202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1204 = 9'he0 == r_count_2_io_out ? io_r_224_b : _GEN_1203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1205 = 9'he1 == r_count_2_io_out ? io_r_225_b : _GEN_1204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1206 = 9'he2 == r_count_2_io_out ? io_r_226_b : _GEN_1205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1207 = 9'he3 == r_count_2_io_out ? io_r_227_b : _GEN_1206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1208 = 9'he4 == r_count_2_io_out ? io_r_228_b : _GEN_1207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1209 = 9'he5 == r_count_2_io_out ? io_r_229_b : _GEN_1208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1210 = 9'he6 == r_count_2_io_out ? io_r_230_b : _GEN_1209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1211 = 9'he7 == r_count_2_io_out ? io_r_231_b : _GEN_1210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1212 = 9'he8 == r_count_2_io_out ? io_r_232_b : _GEN_1211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1213 = 9'he9 == r_count_2_io_out ? io_r_233_b : _GEN_1212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1214 = 9'hea == r_count_2_io_out ? io_r_234_b : _GEN_1213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1215 = 9'heb == r_count_2_io_out ? io_r_235_b : _GEN_1214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1216 = 9'hec == r_count_2_io_out ? io_r_236_b : _GEN_1215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1217 = 9'hed == r_count_2_io_out ? io_r_237_b : _GEN_1216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1218 = 9'hee == r_count_2_io_out ? io_r_238_b : _GEN_1217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1219 = 9'hef == r_count_2_io_out ? io_r_239_b : _GEN_1218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1220 = 9'hf0 == r_count_2_io_out ? io_r_240_b : _GEN_1219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1221 = 9'hf1 == r_count_2_io_out ? io_r_241_b : _GEN_1220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1222 = 9'hf2 == r_count_2_io_out ? io_r_242_b : _GEN_1221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1223 = 9'hf3 == r_count_2_io_out ? io_r_243_b : _GEN_1222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1224 = 9'hf4 == r_count_2_io_out ? io_r_244_b : _GEN_1223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1225 = 9'hf5 == r_count_2_io_out ? io_r_245_b : _GEN_1224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1226 = 9'hf6 == r_count_2_io_out ? io_r_246_b : _GEN_1225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1227 = 9'hf7 == r_count_2_io_out ? io_r_247_b : _GEN_1226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1228 = 9'hf8 == r_count_2_io_out ? io_r_248_b : _GEN_1227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1229 = 9'hf9 == r_count_2_io_out ? io_r_249_b : _GEN_1228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1230 = 9'hfa == r_count_2_io_out ? io_r_250_b : _GEN_1229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1231 = 9'hfb == r_count_2_io_out ? io_r_251_b : _GEN_1230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1232 = 9'hfc == r_count_2_io_out ? io_r_252_b : _GEN_1231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1233 = 9'hfd == r_count_2_io_out ? io_r_253_b : _GEN_1232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1234 = 9'hfe == r_count_2_io_out ? io_r_254_b : _GEN_1233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1235 = 9'hff == r_count_2_io_out ? io_r_255_b : _GEN_1234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1236 = 9'h100 == r_count_2_io_out ? io_r_256_b : _GEN_1235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1237 = 9'h101 == r_count_2_io_out ? io_r_257_b : _GEN_1236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1238 = 9'h102 == r_count_2_io_out ? io_r_258_b : _GEN_1237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1239 = 9'h103 == r_count_2_io_out ? io_r_259_b : _GEN_1238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1240 = 9'h104 == r_count_2_io_out ? io_r_260_b : _GEN_1239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1241 = 9'h105 == r_count_2_io_out ? io_r_261_b : _GEN_1240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1242 = 9'h106 == r_count_2_io_out ? io_r_262_b : _GEN_1241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1243 = 9'h107 == r_count_2_io_out ? io_r_263_b : _GEN_1242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1244 = 9'h108 == r_count_2_io_out ? io_r_264_b : _GEN_1243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1245 = 9'h109 == r_count_2_io_out ? io_r_265_b : _GEN_1244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1246 = 9'h10a == r_count_2_io_out ? io_r_266_b : _GEN_1245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1247 = 9'h10b == r_count_2_io_out ? io_r_267_b : _GEN_1246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1248 = 9'h10c == r_count_2_io_out ? io_r_268_b : _GEN_1247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1249 = 9'h10d == r_count_2_io_out ? io_r_269_b : _GEN_1248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1250 = 9'h10e == r_count_2_io_out ? io_r_270_b : _GEN_1249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1251 = 9'h10f == r_count_2_io_out ? io_r_271_b : _GEN_1250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1252 = 9'h110 == r_count_2_io_out ? io_r_272_b : _GEN_1251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1253 = 9'h111 == r_count_2_io_out ? io_r_273_b : _GEN_1252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1254 = 9'h112 == r_count_2_io_out ? io_r_274_b : _GEN_1253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1255 = 9'h113 == r_count_2_io_out ? io_r_275_b : _GEN_1254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1256 = 9'h114 == r_count_2_io_out ? io_r_276_b : _GEN_1255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1257 = 9'h115 == r_count_2_io_out ? io_r_277_b : _GEN_1256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1258 = 9'h116 == r_count_2_io_out ? io_r_278_b : _GEN_1257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1259 = 9'h117 == r_count_2_io_out ? io_r_279_b : _GEN_1258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1260 = 9'h118 == r_count_2_io_out ? io_r_280_b : _GEN_1259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1261 = 9'h119 == r_count_2_io_out ? io_r_281_b : _GEN_1260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1262 = 9'h11a == r_count_2_io_out ? io_r_282_b : _GEN_1261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1263 = 9'h11b == r_count_2_io_out ? io_r_283_b : _GEN_1262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1264 = 9'h11c == r_count_2_io_out ? io_r_284_b : _GEN_1263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1265 = 9'h11d == r_count_2_io_out ? io_r_285_b : _GEN_1264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1266 = 9'h11e == r_count_2_io_out ? io_r_286_b : _GEN_1265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1267 = 9'h11f == r_count_2_io_out ? io_r_287_b : _GEN_1266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1268 = 9'h120 == r_count_2_io_out ? io_r_288_b : _GEN_1267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1269 = 9'h121 == r_count_2_io_out ? io_r_289_b : _GEN_1268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1270 = 9'h122 == r_count_2_io_out ? io_r_290_b : _GEN_1269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1271 = 9'h123 == r_count_2_io_out ? io_r_291_b : _GEN_1270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1272 = 9'h124 == r_count_2_io_out ? io_r_292_b : _GEN_1271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1273 = 9'h125 == r_count_2_io_out ? io_r_293_b : _GEN_1272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1274 = 9'h126 == r_count_2_io_out ? io_r_294_b : _GEN_1273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1275 = 9'h127 == r_count_2_io_out ? io_r_295_b : _GEN_1274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1276 = 9'h128 == r_count_2_io_out ? io_r_296_b : _GEN_1275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1277 = 9'h129 == r_count_2_io_out ? io_r_297_b : _GEN_1276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1278 = 9'h12a == r_count_2_io_out ? io_r_298_b : _GEN_1277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1279 = 9'h12b == r_count_2_io_out ? io_r_299_b : _GEN_1278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1280 = 9'h12c == r_count_2_io_out ? io_r_300_b : _GEN_1279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1281 = 9'h12d == r_count_2_io_out ? io_r_301_b : _GEN_1280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1282 = 9'h12e == r_count_2_io_out ? io_r_302_b : _GEN_1281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1283 = 9'h12f == r_count_2_io_out ? io_r_303_b : _GEN_1282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1284 = 9'h130 == r_count_2_io_out ? io_r_304_b : _GEN_1283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1285 = 9'h131 == r_count_2_io_out ? io_r_305_b : _GEN_1284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1286 = 9'h132 == r_count_2_io_out ? io_r_306_b : _GEN_1285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1287 = 9'h133 == r_count_2_io_out ? io_r_307_b : _GEN_1286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1288 = 9'h134 == r_count_2_io_out ? io_r_308_b : _GEN_1287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1289 = 9'h135 == r_count_2_io_out ? io_r_309_b : _GEN_1288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1290 = 9'h136 == r_count_2_io_out ? io_r_310_b : _GEN_1289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1291 = 9'h137 == r_count_2_io_out ? io_r_311_b : _GEN_1290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1292 = 9'h138 == r_count_2_io_out ? io_r_312_b : _GEN_1291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1293 = 9'h139 == r_count_2_io_out ? io_r_313_b : _GEN_1292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1294 = 9'h13a == r_count_2_io_out ? io_r_314_b : _GEN_1293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1295 = 9'h13b == r_count_2_io_out ? io_r_315_b : _GEN_1294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1296 = 9'h13c == r_count_2_io_out ? io_r_316_b : _GEN_1295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1297 = 9'h13d == r_count_2_io_out ? io_r_317_b : _GEN_1296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1298 = 9'h13e == r_count_2_io_out ? io_r_318_b : _GEN_1297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1299 = 9'h13f == r_count_2_io_out ? io_r_319_b : _GEN_1298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1300 = 9'h140 == r_count_2_io_out ? io_r_320_b : _GEN_1299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1301 = 9'h141 == r_count_2_io_out ? io_r_321_b : _GEN_1300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1302 = 9'h142 == r_count_2_io_out ? io_r_322_b : _GEN_1301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1303 = 9'h143 == r_count_2_io_out ? io_r_323_b : _GEN_1302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1304 = 9'h144 == r_count_2_io_out ? io_r_324_b : _GEN_1303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1305 = 9'h145 == r_count_2_io_out ? io_r_325_b : _GEN_1304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1306 = 9'h146 == r_count_2_io_out ? io_r_326_b : _GEN_1305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1307 = 9'h147 == r_count_2_io_out ? io_r_327_b : _GEN_1306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1308 = 9'h148 == r_count_2_io_out ? io_r_328_b : _GEN_1307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1309 = 9'h149 == r_count_2_io_out ? io_r_329_b : _GEN_1308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1310 = 9'h14a == r_count_2_io_out ? io_r_330_b : _GEN_1309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1311 = 9'h14b == r_count_2_io_out ? io_r_331_b : _GEN_1310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1312 = 9'h14c == r_count_2_io_out ? io_r_332_b : _GEN_1311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1313 = 9'h14d == r_count_2_io_out ? io_r_333_b : _GEN_1312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1314 = 9'h14e == r_count_2_io_out ? io_r_334_b : _GEN_1313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1315 = 9'h14f == r_count_2_io_out ? io_r_335_b : _GEN_1314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1316 = 9'h150 == r_count_2_io_out ? io_r_336_b : _GEN_1315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1317 = 9'h151 == r_count_2_io_out ? io_r_337_b : _GEN_1316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1318 = 9'h152 == r_count_2_io_out ? io_r_338_b : _GEN_1317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1319 = 9'h153 == r_count_2_io_out ? io_r_339_b : _GEN_1318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1320 = 9'h154 == r_count_2_io_out ? io_r_340_b : _GEN_1319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1321 = 9'h155 == r_count_2_io_out ? io_r_341_b : _GEN_1320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1322 = 9'h156 == r_count_2_io_out ? io_r_342_b : _GEN_1321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1323 = 9'h157 == r_count_2_io_out ? io_r_343_b : _GEN_1322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1324 = 9'h158 == r_count_2_io_out ? io_r_344_b : _GEN_1323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1325 = 9'h159 == r_count_2_io_out ? io_r_345_b : _GEN_1324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1326 = 9'h15a == r_count_2_io_out ? io_r_346_b : _GEN_1325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1327 = 9'h15b == r_count_2_io_out ? io_r_347_b : _GEN_1326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1328 = 9'h15c == r_count_2_io_out ? io_r_348_b : _GEN_1327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1329 = 9'h15d == r_count_2_io_out ? io_r_349_b : _GEN_1328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1330 = 9'h15e == r_count_2_io_out ? io_r_350_b : _GEN_1329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1331 = 9'h15f == r_count_2_io_out ? io_r_351_b : _GEN_1330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1332 = 9'h160 == r_count_2_io_out ? io_r_352_b : _GEN_1331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1333 = 9'h161 == r_count_2_io_out ? io_r_353_b : _GEN_1332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1334 = 9'h162 == r_count_2_io_out ? io_r_354_b : _GEN_1333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1335 = 9'h163 == r_count_2_io_out ? io_r_355_b : _GEN_1334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1336 = 9'h164 == r_count_2_io_out ? io_r_356_b : _GEN_1335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1337 = 9'h165 == r_count_2_io_out ? io_r_357_b : _GEN_1336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1338 = 9'h166 == r_count_2_io_out ? io_r_358_b : _GEN_1337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1339 = 9'h167 == r_count_2_io_out ? io_r_359_b : _GEN_1338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1340 = 9'h168 == r_count_2_io_out ? io_r_360_b : _GEN_1339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1341 = 9'h169 == r_count_2_io_out ? io_r_361_b : _GEN_1340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1342 = 9'h16a == r_count_2_io_out ? io_r_362_b : _GEN_1341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1343 = 9'h16b == r_count_2_io_out ? io_r_363_b : _GEN_1342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1344 = 9'h16c == r_count_2_io_out ? io_r_364_b : _GEN_1343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1345 = 9'h16d == r_count_2_io_out ? io_r_365_b : _GEN_1344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1346 = 9'h16e == r_count_2_io_out ? io_r_366_b : _GEN_1345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1347 = 9'h16f == r_count_2_io_out ? io_r_367_b : _GEN_1346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1348 = 9'h170 == r_count_2_io_out ? io_r_368_b : _GEN_1347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1349 = 9'h171 == r_count_2_io_out ? io_r_369_b : _GEN_1348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1350 = 9'h172 == r_count_2_io_out ? io_r_370_b : _GEN_1349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1351 = 9'h173 == r_count_2_io_out ? io_r_371_b : _GEN_1350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1352 = 9'h174 == r_count_2_io_out ? io_r_372_b : _GEN_1351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1353 = 9'h175 == r_count_2_io_out ? io_r_373_b : _GEN_1352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1354 = 9'h176 == r_count_2_io_out ? io_r_374_b : _GEN_1353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1355 = 9'h177 == r_count_2_io_out ? io_r_375_b : _GEN_1354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1356 = 9'h178 == r_count_2_io_out ? io_r_376_b : _GEN_1355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1357 = 9'h179 == r_count_2_io_out ? io_r_377_b : _GEN_1356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1358 = 9'h17a == r_count_2_io_out ? io_r_378_b : _GEN_1357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1359 = 9'h17b == r_count_2_io_out ? io_r_379_b : _GEN_1358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1360 = 9'h17c == r_count_2_io_out ? io_r_380_b : _GEN_1359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1361 = 9'h17d == r_count_2_io_out ? io_r_381_b : _GEN_1360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1362 = 9'h17e == r_count_2_io_out ? io_r_382_b : _GEN_1361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1363 = 9'h17f == r_count_2_io_out ? io_r_383_b : _GEN_1362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1364 = 9'h180 == r_count_2_io_out ? io_r_384_b : _GEN_1363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1365 = 9'h181 == r_count_2_io_out ? io_r_385_b : _GEN_1364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1366 = 9'h182 == r_count_2_io_out ? io_r_386_b : _GEN_1365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1367 = 9'h183 == r_count_2_io_out ? io_r_387_b : _GEN_1366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1368 = 9'h184 == r_count_2_io_out ? io_r_388_b : _GEN_1367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1369 = 9'h185 == r_count_2_io_out ? io_r_389_b : _GEN_1368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1370 = 9'h186 == r_count_2_io_out ? io_r_390_b : _GEN_1369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1371 = 9'h187 == r_count_2_io_out ? io_r_391_b : _GEN_1370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1372 = 9'h188 == r_count_2_io_out ? io_r_392_b : _GEN_1371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1373 = 9'h189 == r_count_2_io_out ? io_r_393_b : _GEN_1372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1374 = 9'h18a == r_count_2_io_out ? io_r_394_b : _GEN_1373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1375 = 9'h18b == r_count_2_io_out ? io_r_395_b : _GEN_1374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1376 = 9'h18c == r_count_2_io_out ? io_r_396_b : _GEN_1375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1377 = 9'h18d == r_count_2_io_out ? io_r_397_b : _GEN_1376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1378 = 9'h18e == r_count_2_io_out ? io_r_398_b : _GEN_1377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1381 = 9'h1 == r_count_3_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1382 = 9'h2 == r_count_3_io_out ? io_r_2_b : _GEN_1381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1383 = 9'h3 == r_count_3_io_out ? io_r_3_b : _GEN_1382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1384 = 9'h4 == r_count_3_io_out ? io_r_4_b : _GEN_1383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1385 = 9'h5 == r_count_3_io_out ? io_r_5_b : _GEN_1384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1386 = 9'h6 == r_count_3_io_out ? io_r_6_b : _GEN_1385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1387 = 9'h7 == r_count_3_io_out ? io_r_7_b : _GEN_1386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1388 = 9'h8 == r_count_3_io_out ? io_r_8_b : _GEN_1387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1389 = 9'h9 == r_count_3_io_out ? io_r_9_b : _GEN_1388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1390 = 9'ha == r_count_3_io_out ? io_r_10_b : _GEN_1389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1391 = 9'hb == r_count_3_io_out ? io_r_11_b : _GEN_1390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1392 = 9'hc == r_count_3_io_out ? io_r_12_b : _GEN_1391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1393 = 9'hd == r_count_3_io_out ? io_r_13_b : _GEN_1392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1394 = 9'he == r_count_3_io_out ? io_r_14_b : _GEN_1393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1395 = 9'hf == r_count_3_io_out ? io_r_15_b : _GEN_1394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1396 = 9'h10 == r_count_3_io_out ? io_r_16_b : _GEN_1395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1397 = 9'h11 == r_count_3_io_out ? io_r_17_b : _GEN_1396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1398 = 9'h12 == r_count_3_io_out ? io_r_18_b : _GEN_1397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1399 = 9'h13 == r_count_3_io_out ? io_r_19_b : _GEN_1398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1400 = 9'h14 == r_count_3_io_out ? io_r_20_b : _GEN_1399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1401 = 9'h15 == r_count_3_io_out ? io_r_21_b : _GEN_1400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1402 = 9'h16 == r_count_3_io_out ? io_r_22_b : _GEN_1401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1403 = 9'h17 == r_count_3_io_out ? io_r_23_b : _GEN_1402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1404 = 9'h18 == r_count_3_io_out ? io_r_24_b : _GEN_1403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1405 = 9'h19 == r_count_3_io_out ? io_r_25_b : _GEN_1404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1406 = 9'h1a == r_count_3_io_out ? io_r_26_b : _GEN_1405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1407 = 9'h1b == r_count_3_io_out ? io_r_27_b : _GEN_1406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1408 = 9'h1c == r_count_3_io_out ? io_r_28_b : _GEN_1407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1409 = 9'h1d == r_count_3_io_out ? io_r_29_b : _GEN_1408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1410 = 9'h1e == r_count_3_io_out ? io_r_30_b : _GEN_1409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1411 = 9'h1f == r_count_3_io_out ? io_r_31_b : _GEN_1410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1412 = 9'h20 == r_count_3_io_out ? io_r_32_b : _GEN_1411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1413 = 9'h21 == r_count_3_io_out ? io_r_33_b : _GEN_1412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1414 = 9'h22 == r_count_3_io_out ? io_r_34_b : _GEN_1413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1415 = 9'h23 == r_count_3_io_out ? io_r_35_b : _GEN_1414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1416 = 9'h24 == r_count_3_io_out ? io_r_36_b : _GEN_1415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1417 = 9'h25 == r_count_3_io_out ? io_r_37_b : _GEN_1416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1418 = 9'h26 == r_count_3_io_out ? io_r_38_b : _GEN_1417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1419 = 9'h27 == r_count_3_io_out ? io_r_39_b : _GEN_1418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1420 = 9'h28 == r_count_3_io_out ? io_r_40_b : _GEN_1419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1421 = 9'h29 == r_count_3_io_out ? io_r_41_b : _GEN_1420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1422 = 9'h2a == r_count_3_io_out ? io_r_42_b : _GEN_1421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1423 = 9'h2b == r_count_3_io_out ? io_r_43_b : _GEN_1422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1424 = 9'h2c == r_count_3_io_out ? io_r_44_b : _GEN_1423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1425 = 9'h2d == r_count_3_io_out ? io_r_45_b : _GEN_1424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1426 = 9'h2e == r_count_3_io_out ? io_r_46_b : _GEN_1425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1427 = 9'h2f == r_count_3_io_out ? io_r_47_b : _GEN_1426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1428 = 9'h30 == r_count_3_io_out ? io_r_48_b : _GEN_1427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1429 = 9'h31 == r_count_3_io_out ? io_r_49_b : _GEN_1428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1430 = 9'h32 == r_count_3_io_out ? io_r_50_b : _GEN_1429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1431 = 9'h33 == r_count_3_io_out ? io_r_51_b : _GEN_1430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1432 = 9'h34 == r_count_3_io_out ? io_r_52_b : _GEN_1431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1433 = 9'h35 == r_count_3_io_out ? io_r_53_b : _GEN_1432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1434 = 9'h36 == r_count_3_io_out ? io_r_54_b : _GEN_1433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1435 = 9'h37 == r_count_3_io_out ? io_r_55_b : _GEN_1434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1436 = 9'h38 == r_count_3_io_out ? io_r_56_b : _GEN_1435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1437 = 9'h39 == r_count_3_io_out ? io_r_57_b : _GEN_1436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1438 = 9'h3a == r_count_3_io_out ? io_r_58_b : _GEN_1437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1439 = 9'h3b == r_count_3_io_out ? io_r_59_b : _GEN_1438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1440 = 9'h3c == r_count_3_io_out ? io_r_60_b : _GEN_1439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1441 = 9'h3d == r_count_3_io_out ? io_r_61_b : _GEN_1440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1442 = 9'h3e == r_count_3_io_out ? io_r_62_b : _GEN_1441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1443 = 9'h3f == r_count_3_io_out ? io_r_63_b : _GEN_1442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1444 = 9'h40 == r_count_3_io_out ? io_r_64_b : _GEN_1443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1445 = 9'h41 == r_count_3_io_out ? io_r_65_b : _GEN_1444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1446 = 9'h42 == r_count_3_io_out ? io_r_66_b : _GEN_1445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1447 = 9'h43 == r_count_3_io_out ? io_r_67_b : _GEN_1446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1448 = 9'h44 == r_count_3_io_out ? io_r_68_b : _GEN_1447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1449 = 9'h45 == r_count_3_io_out ? io_r_69_b : _GEN_1448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1450 = 9'h46 == r_count_3_io_out ? io_r_70_b : _GEN_1449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1451 = 9'h47 == r_count_3_io_out ? io_r_71_b : _GEN_1450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1452 = 9'h48 == r_count_3_io_out ? io_r_72_b : _GEN_1451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1453 = 9'h49 == r_count_3_io_out ? io_r_73_b : _GEN_1452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1454 = 9'h4a == r_count_3_io_out ? io_r_74_b : _GEN_1453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1455 = 9'h4b == r_count_3_io_out ? io_r_75_b : _GEN_1454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1456 = 9'h4c == r_count_3_io_out ? io_r_76_b : _GEN_1455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1457 = 9'h4d == r_count_3_io_out ? io_r_77_b : _GEN_1456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1458 = 9'h4e == r_count_3_io_out ? io_r_78_b : _GEN_1457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1459 = 9'h4f == r_count_3_io_out ? io_r_79_b : _GEN_1458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1460 = 9'h50 == r_count_3_io_out ? io_r_80_b : _GEN_1459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1461 = 9'h51 == r_count_3_io_out ? io_r_81_b : _GEN_1460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1462 = 9'h52 == r_count_3_io_out ? io_r_82_b : _GEN_1461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1463 = 9'h53 == r_count_3_io_out ? io_r_83_b : _GEN_1462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1464 = 9'h54 == r_count_3_io_out ? io_r_84_b : _GEN_1463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1465 = 9'h55 == r_count_3_io_out ? io_r_85_b : _GEN_1464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1466 = 9'h56 == r_count_3_io_out ? io_r_86_b : _GEN_1465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1467 = 9'h57 == r_count_3_io_out ? io_r_87_b : _GEN_1466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1468 = 9'h58 == r_count_3_io_out ? io_r_88_b : _GEN_1467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1469 = 9'h59 == r_count_3_io_out ? io_r_89_b : _GEN_1468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1470 = 9'h5a == r_count_3_io_out ? io_r_90_b : _GEN_1469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1471 = 9'h5b == r_count_3_io_out ? io_r_91_b : _GEN_1470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1472 = 9'h5c == r_count_3_io_out ? io_r_92_b : _GEN_1471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1473 = 9'h5d == r_count_3_io_out ? io_r_93_b : _GEN_1472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1474 = 9'h5e == r_count_3_io_out ? io_r_94_b : _GEN_1473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1475 = 9'h5f == r_count_3_io_out ? io_r_95_b : _GEN_1474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1476 = 9'h60 == r_count_3_io_out ? io_r_96_b : _GEN_1475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1477 = 9'h61 == r_count_3_io_out ? io_r_97_b : _GEN_1476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1478 = 9'h62 == r_count_3_io_out ? io_r_98_b : _GEN_1477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1479 = 9'h63 == r_count_3_io_out ? io_r_99_b : _GEN_1478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1480 = 9'h64 == r_count_3_io_out ? io_r_100_b : _GEN_1479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1481 = 9'h65 == r_count_3_io_out ? io_r_101_b : _GEN_1480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1482 = 9'h66 == r_count_3_io_out ? io_r_102_b : _GEN_1481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1483 = 9'h67 == r_count_3_io_out ? io_r_103_b : _GEN_1482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1484 = 9'h68 == r_count_3_io_out ? io_r_104_b : _GEN_1483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1485 = 9'h69 == r_count_3_io_out ? io_r_105_b : _GEN_1484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1486 = 9'h6a == r_count_3_io_out ? io_r_106_b : _GEN_1485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1487 = 9'h6b == r_count_3_io_out ? io_r_107_b : _GEN_1486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1488 = 9'h6c == r_count_3_io_out ? io_r_108_b : _GEN_1487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1489 = 9'h6d == r_count_3_io_out ? io_r_109_b : _GEN_1488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1490 = 9'h6e == r_count_3_io_out ? io_r_110_b : _GEN_1489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1491 = 9'h6f == r_count_3_io_out ? io_r_111_b : _GEN_1490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1492 = 9'h70 == r_count_3_io_out ? io_r_112_b : _GEN_1491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1493 = 9'h71 == r_count_3_io_out ? io_r_113_b : _GEN_1492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1494 = 9'h72 == r_count_3_io_out ? io_r_114_b : _GEN_1493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1495 = 9'h73 == r_count_3_io_out ? io_r_115_b : _GEN_1494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1496 = 9'h74 == r_count_3_io_out ? io_r_116_b : _GEN_1495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1497 = 9'h75 == r_count_3_io_out ? io_r_117_b : _GEN_1496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1498 = 9'h76 == r_count_3_io_out ? io_r_118_b : _GEN_1497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1499 = 9'h77 == r_count_3_io_out ? io_r_119_b : _GEN_1498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1500 = 9'h78 == r_count_3_io_out ? io_r_120_b : _GEN_1499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1501 = 9'h79 == r_count_3_io_out ? io_r_121_b : _GEN_1500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1502 = 9'h7a == r_count_3_io_out ? io_r_122_b : _GEN_1501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1503 = 9'h7b == r_count_3_io_out ? io_r_123_b : _GEN_1502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1504 = 9'h7c == r_count_3_io_out ? io_r_124_b : _GEN_1503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1505 = 9'h7d == r_count_3_io_out ? io_r_125_b : _GEN_1504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1506 = 9'h7e == r_count_3_io_out ? io_r_126_b : _GEN_1505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1507 = 9'h7f == r_count_3_io_out ? io_r_127_b : _GEN_1506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1508 = 9'h80 == r_count_3_io_out ? io_r_128_b : _GEN_1507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1509 = 9'h81 == r_count_3_io_out ? io_r_129_b : _GEN_1508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1510 = 9'h82 == r_count_3_io_out ? io_r_130_b : _GEN_1509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1511 = 9'h83 == r_count_3_io_out ? io_r_131_b : _GEN_1510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1512 = 9'h84 == r_count_3_io_out ? io_r_132_b : _GEN_1511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1513 = 9'h85 == r_count_3_io_out ? io_r_133_b : _GEN_1512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1514 = 9'h86 == r_count_3_io_out ? io_r_134_b : _GEN_1513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1515 = 9'h87 == r_count_3_io_out ? io_r_135_b : _GEN_1514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1516 = 9'h88 == r_count_3_io_out ? io_r_136_b : _GEN_1515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1517 = 9'h89 == r_count_3_io_out ? io_r_137_b : _GEN_1516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1518 = 9'h8a == r_count_3_io_out ? io_r_138_b : _GEN_1517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1519 = 9'h8b == r_count_3_io_out ? io_r_139_b : _GEN_1518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1520 = 9'h8c == r_count_3_io_out ? io_r_140_b : _GEN_1519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1521 = 9'h8d == r_count_3_io_out ? io_r_141_b : _GEN_1520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1522 = 9'h8e == r_count_3_io_out ? io_r_142_b : _GEN_1521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1523 = 9'h8f == r_count_3_io_out ? io_r_143_b : _GEN_1522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1524 = 9'h90 == r_count_3_io_out ? io_r_144_b : _GEN_1523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1525 = 9'h91 == r_count_3_io_out ? io_r_145_b : _GEN_1524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1526 = 9'h92 == r_count_3_io_out ? io_r_146_b : _GEN_1525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1527 = 9'h93 == r_count_3_io_out ? io_r_147_b : _GEN_1526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1528 = 9'h94 == r_count_3_io_out ? io_r_148_b : _GEN_1527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1529 = 9'h95 == r_count_3_io_out ? io_r_149_b : _GEN_1528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1530 = 9'h96 == r_count_3_io_out ? io_r_150_b : _GEN_1529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1531 = 9'h97 == r_count_3_io_out ? io_r_151_b : _GEN_1530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1532 = 9'h98 == r_count_3_io_out ? io_r_152_b : _GEN_1531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1533 = 9'h99 == r_count_3_io_out ? io_r_153_b : _GEN_1532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1534 = 9'h9a == r_count_3_io_out ? io_r_154_b : _GEN_1533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1535 = 9'h9b == r_count_3_io_out ? io_r_155_b : _GEN_1534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1536 = 9'h9c == r_count_3_io_out ? io_r_156_b : _GEN_1535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1537 = 9'h9d == r_count_3_io_out ? io_r_157_b : _GEN_1536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1538 = 9'h9e == r_count_3_io_out ? io_r_158_b : _GEN_1537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1539 = 9'h9f == r_count_3_io_out ? io_r_159_b : _GEN_1538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1540 = 9'ha0 == r_count_3_io_out ? io_r_160_b : _GEN_1539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1541 = 9'ha1 == r_count_3_io_out ? io_r_161_b : _GEN_1540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1542 = 9'ha2 == r_count_3_io_out ? io_r_162_b : _GEN_1541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1543 = 9'ha3 == r_count_3_io_out ? io_r_163_b : _GEN_1542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1544 = 9'ha4 == r_count_3_io_out ? io_r_164_b : _GEN_1543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1545 = 9'ha5 == r_count_3_io_out ? io_r_165_b : _GEN_1544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1546 = 9'ha6 == r_count_3_io_out ? io_r_166_b : _GEN_1545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1547 = 9'ha7 == r_count_3_io_out ? io_r_167_b : _GEN_1546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1548 = 9'ha8 == r_count_3_io_out ? io_r_168_b : _GEN_1547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1549 = 9'ha9 == r_count_3_io_out ? io_r_169_b : _GEN_1548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1550 = 9'haa == r_count_3_io_out ? io_r_170_b : _GEN_1549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1551 = 9'hab == r_count_3_io_out ? io_r_171_b : _GEN_1550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1552 = 9'hac == r_count_3_io_out ? io_r_172_b : _GEN_1551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1553 = 9'had == r_count_3_io_out ? io_r_173_b : _GEN_1552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1554 = 9'hae == r_count_3_io_out ? io_r_174_b : _GEN_1553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1555 = 9'haf == r_count_3_io_out ? io_r_175_b : _GEN_1554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1556 = 9'hb0 == r_count_3_io_out ? io_r_176_b : _GEN_1555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1557 = 9'hb1 == r_count_3_io_out ? io_r_177_b : _GEN_1556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1558 = 9'hb2 == r_count_3_io_out ? io_r_178_b : _GEN_1557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1559 = 9'hb3 == r_count_3_io_out ? io_r_179_b : _GEN_1558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1560 = 9'hb4 == r_count_3_io_out ? io_r_180_b : _GEN_1559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1561 = 9'hb5 == r_count_3_io_out ? io_r_181_b : _GEN_1560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1562 = 9'hb6 == r_count_3_io_out ? io_r_182_b : _GEN_1561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1563 = 9'hb7 == r_count_3_io_out ? io_r_183_b : _GEN_1562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1564 = 9'hb8 == r_count_3_io_out ? io_r_184_b : _GEN_1563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1565 = 9'hb9 == r_count_3_io_out ? io_r_185_b : _GEN_1564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1566 = 9'hba == r_count_3_io_out ? io_r_186_b : _GEN_1565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1567 = 9'hbb == r_count_3_io_out ? io_r_187_b : _GEN_1566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1568 = 9'hbc == r_count_3_io_out ? io_r_188_b : _GEN_1567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1569 = 9'hbd == r_count_3_io_out ? io_r_189_b : _GEN_1568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1570 = 9'hbe == r_count_3_io_out ? io_r_190_b : _GEN_1569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1571 = 9'hbf == r_count_3_io_out ? io_r_191_b : _GEN_1570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1572 = 9'hc0 == r_count_3_io_out ? io_r_192_b : _GEN_1571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1573 = 9'hc1 == r_count_3_io_out ? io_r_193_b : _GEN_1572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1574 = 9'hc2 == r_count_3_io_out ? io_r_194_b : _GEN_1573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1575 = 9'hc3 == r_count_3_io_out ? io_r_195_b : _GEN_1574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1576 = 9'hc4 == r_count_3_io_out ? io_r_196_b : _GEN_1575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1577 = 9'hc5 == r_count_3_io_out ? io_r_197_b : _GEN_1576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1578 = 9'hc6 == r_count_3_io_out ? io_r_198_b : _GEN_1577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1579 = 9'hc7 == r_count_3_io_out ? io_r_199_b : _GEN_1578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1580 = 9'hc8 == r_count_3_io_out ? io_r_200_b : _GEN_1579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1581 = 9'hc9 == r_count_3_io_out ? io_r_201_b : _GEN_1580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1582 = 9'hca == r_count_3_io_out ? io_r_202_b : _GEN_1581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1583 = 9'hcb == r_count_3_io_out ? io_r_203_b : _GEN_1582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1584 = 9'hcc == r_count_3_io_out ? io_r_204_b : _GEN_1583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1585 = 9'hcd == r_count_3_io_out ? io_r_205_b : _GEN_1584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1586 = 9'hce == r_count_3_io_out ? io_r_206_b : _GEN_1585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1587 = 9'hcf == r_count_3_io_out ? io_r_207_b : _GEN_1586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1588 = 9'hd0 == r_count_3_io_out ? io_r_208_b : _GEN_1587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1589 = 9'hd1 == r_count_3_io_out ? io_r_209_b : _GEN_1588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1590 = 9'hd2 == r_count_3_io_out ? io_r_210_b : _GEN_1589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1591 = 9'hd3 == r_count_3_io_out ? io_r_211_b : _GEN_1590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1592 = 9'hd4 == r_count_3_io_out ? io_r_212_b : _GEN_1591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1593 = 9'hd5 == r_count_3_io_out ? io_r_213_b : _GEN_1592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1594 = 9'hd6 == r_count_3_io_out ? io_r_214_b : _GEN_1593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1595 = 9'hd7 == r_count_3_io_out ? io_r_215_b : _GEN_1594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1596 = 9'hd8 == r_count_3_io_out ? io_r_216_b : _GEN_1595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1597 = 9'hd9 == r_count_3_io_out ? io_r_217_b : _GEN_1596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1598 = 9'hda == r_count_3_io_out ? io_r_218_b : _GEN_1597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1599 = 9'hdb == r_count_3_io_out ? io_r_219_b : _GEN_1598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1600 = 9'hdc == r_count_3_io_out ? io_r_220_b : _GEN_1599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1601 = 9'hdd == r_count_3_io_out ? io_r_221_b : _GEN_1600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1602 = 9'hde == r_count_3_io_out ? io_r_222_b : _GEN_1601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1603 = 9'hdf == r_count_3_io_out ? io_r_223_b : _GEN_1602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1604 = 9'he0 == r_count_3_io_out ? io_r_224_b : _GEN_1603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1605 = 9'he1 == r_count_3_io_out ? io_r_225_b : _GEN_1604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1606 = 9'he2 == r_count_3_io_out ? io_r_226_b : _GEN_1605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1607 = 9'he3 == r_count_3_io_out ? io_r_227_b : _GEN_1606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1608 = 9'he4 == r_count_3_io_out ? io_r_228_b : _GEN_1607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1609 = 9'he5 == r_count_3_io_out ? io_r_229_b : _GEN_1608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1610 = 9'he6 == r_count_3_io_out ? io_r_230_b : _GEN_1609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1611 = 9'he7 == r_count_3_io_out ? io_r_231_b : _GEN_1610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1612 = 9'he8 == r_count_3_io_out ? io_r_232_b : _GEN_1611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1613 = 9'he9 == r_count_3_io_out ? io_r_233_b : _GEN_1612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1614 = 9'hea == r_count_3_io_out ? io_r_234_b : _GEN_1613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1615 = 9'heb == r_count_3_io_out ? io_r_235_b : _GEN_1614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1616 = 9'hec == r_count_3_io_out ? io_r_236_b : _GEN_1615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1617 = 9'hed == r_count_3_io_out ? io_r_237_b : _GEN_1616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1618 = 9'hee == r_count_3_io_out ? io_r_238_b : _GEN_1617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1619 = 9'hef == r_count_3_io_out ? io_r_239_b : _GEN_1618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1620 = 9'hf0 == r_count_3_io_out ? io_r_240_b : _GEN_1619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1621 = 9'hf1 == r_count_3_io_out ? io_r_241_b : _GEN_1620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1622 = 9'hf2 == r_count_3_io_out ? io_r_242_b : _GEN_1621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1623 = 9'hf3 == r_count_3_io_out ? io_r_243_b : _GEN_1622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1624 = 9'hf4 == r_count_3_io_out ? io_r_244_b : _GEN_1623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1625 = 9'hf5 == r_count_3_io_out ? io_r_245_b : _GEN_1624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1626 = 9'hf6 == r_count_3_io_out ? io_r_246_b : _GEN_1625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1627 = 9'hf7 == r_count_3_io_out ? io_r_247_b : _GEN_1626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1628 = 9'hf8 == r_count_3_io_out ? io_r_248_b : _GEN_1627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1629 = 9'hf9 == r_count_3_io_out ? io_r_249_b : _GEN_1628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1630 = 9'hfa == r_count_3_io_out ? io_r_250_b : _GEN_1629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1631 = 9'hfb == r_count_3_io_out ? io_r_251_b : _GEN_1630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1632 = 9'hfc == r_count_3_io_out ? io_r_252_b : _GEN_1631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1633 = 9'hfd == r_count_3_io_out ? io_r_253_b : _GEN_1632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1634 = 9'hfe == r_count_3_io_out ? io_r_254_b : _GEN_1633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1635 = 9'hff == r_count_3_io_out ? io_r_255_b : _GEN_1634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1636 = 9'h100 == r_count_3_io_out ? io_r_256_b : _GEN_1635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1637 = 9'h101 == r_count_3_io_out ? io_r_257_b : _GEN_1636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1638 = 9'h102 == r_count_3_io_out ? io_r_258_b : _GEN_1637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1639 = 9'h103 == r_count_3_io_out ? io_r_259_b : _GEN_1638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1640 = 9'h104 == r_count_3_io_out ? io_r_260_b : _GEN_1639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1641 = 9'h105 == r_count_3_io_out ? io_r_261_b : _GEN_1640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1642 = 9'h106 == r_count_3_io_out ? io_r_262_b : _GEN_1641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1643 = 9'h107 == r_count_3_io_out ? io_r_263_b : _GEN_1642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1644 = 9'h108 == r_count_3_io_out ? io_r_264_b : _GEN_1643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1645 = 9'h109 == r_count_3_io_out ? io_r_265_b : _GEN_1644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1646 = 9'h10a == r_count_3_io_out ? io_r_266_b : _GEN_1645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1647 = 9'h10b == r_count_3_io_out ? io_r_267_b : _GEN_1646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1648 = 9'h10c == r_count_3_io_out ? io_r_268_b : _GEN_1647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1649 = 9'h10d == r_count_3_io_out ? io_r_269_b : _GEN_1648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1650 = 9'h10e == r_count_3_io_out ? io_r_270_b : _GEN_1649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1651 = 9'h10f == r_count_3_io_out ? io_r_271_b : _GEN_1650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1652 = 9'h110 == r_count_3_io_out ? io_r_272_b : _GEN_1651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1653 = 9'h111 == r_count_3_io_out ? io_r_273_b : _GEN_1652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1654 = 9'h112 == r_count_3_io_out ? io_r_274_b : _GEN_1653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1655 = 9'h113 == r_count_3_io_out ? io_r_275_b : _GEN_1654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1656 = 9'h114 == r_count_3_io_out ? io_r_276_b : _GEN_1655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1657 = 9'h115 == r_count_3_io_out ? io_r_277_b : _GEN_1656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1658 = 9'h116 == r_count_3_io_out ? io_r_278_b : _GEN_1657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1659 = 9'h117 == r_count_3_io_out ? io_r_279_b : _GEN_1658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1660 = 9'h118 == r_count_3_io_out ? io_r_280_b : _GEN_1659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1661 = 9'h119 == r_count_3_io_out ? io_r_281_b : _GEN_1660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1662 = 9'h11a == r_count_3_io_out ? io_r_282_b : _GEN_1661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1663 = 9'h11b == r_count_3_io_out ? io_r_283_b : _GEN_1662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1664 = 9'h11c == r_count_3_io_out ? io_r_284_b : _GEN_1663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1665 = 9'h11d == r_count_3_io_out ? io_r_285_b : _GEN_1664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1666 = 9'h11e == r_count_3_io_out ? io_r_286_b : _GEN_1665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1667 = 9'h11f == r_count_3_io_out ? io_r_287_b : _GEN_1666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1668 = 9'h120 == r_count_3_io_out ? io_r_288_b : _GEN_1667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1669 = 9'h121 == r_count_3_io_out ? io_r_289_b : _GEN_1668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1670 = 9'h122 == r_count_3_io_out ? io_r_290_b : _GEN_1669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1671 = 9'h123 == r_count_3_io_out ? io_r_291_b : _GEN_1670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1672 = 9'h124 == r_count_3_io_out ? io_r_292_b : _GEN_1671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1673 = 9'h125 == r_count_3_io_out ? io_r_293_b : _GEN_1672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1674 = 9'h126 == r_count_3_io_out ? io_r_294_b : _GEN_1673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1675 = 9'h127 == r_count_3_io_out ? io_r_295_b : _GEN_1674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1676 = 9'h128 == r_count_3_io_out ? io_r_296_b : _GEN_1675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1677 = 9'h129 == r_count_3_io_out ? io_r_297_b : _GEN_1676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1678 = 9'h12a == r_count_3_io_out ? io_r_298_b : _GEN_1677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1679 = 9'h12b == r_count_3_io_out ? io_r_299_b : _GEN_1678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1680 = 9'h12c == r_count_3_io_out ? io_r_300_b : _GEN_1679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1681 = 9'h12d == r_count_3_io_out ? io_r_301_b : _GEN_1680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1682 = 9'h12e == r_count_3_io_out ? io_r_302_b : _GEN_1681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1683 = 9'h12f == r_count_3_io_out ? io_r_303_b : _GEN_1682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1684 = 9'h130 == r_count_3_io_out ? io_r_304_b : _GEN_1683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1685 = 9'h131 == r_count_3_io_out ? io_r_305_b : _GEN_1684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1686 = 9'h132 == r_count_3_io_out ? io_r_306_b : _GEN_1685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1687 = 9'h133 == r_count_3_io_out ? io_r_307_b : _GEN_1686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1688 = 9'h134 == r_count_3_io_out ? io_r_308_b : _GEN_1687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1689 = 9'h135 == r_count_3_io_out ? io_r_309_b : _GEN_1688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1690 = 9'h136 == r_count_3_io_out ? io_r_310_b : _GEN_1689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1691 = 9'h137 == r_count_3_io_out ? io_r_311_b : _GEN_1690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1692 = 9'h138 == r_count_3_io_out ? io_r_312_b : _GEN_1691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1693 = 9'h139 == r_count_3_io_out ? io_r_313_b : _GEN_1692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1694 = 9'h13a == r_count_3_io_out ? io_r_314_b : _GEN_1693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1695 = 9'h13b == r_count_3_io_out ? io_r_315_b : _GEN_1694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1696 = 9'h13c == r_count_3_io_out ? io_r_316_b : _GEN_1695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1697 = 9'h13d == r_count_3_io_out ? io_r_317_b : _GEN_1696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1698 = 9'h13e == r_count_3_io_out ? io_r_318_b : _GEN_1697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1699 = 9'h13f == r_count_3_io_out ? io_r_319_b : _GEN_1698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1700 = 9'h140 == r_count_3_io_out ? io_r_320_b : _GEN_1699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1701 = 9'h141 == r_count_3_io_out ? io_r_321_b : _GEN_1700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1702 = 9'h142 == r_count_3_io_out ? io_r_322_b : _GEN_1701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1703 = 9'h143 == r_count_3_io_out ? io_r_323_b : _GEN_1702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1704 = 9'h144 == r_count_3_io_out ? io_r_324_b : _GEN_1703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1705 = 9'h145 == r_count_3_io_out ? io_r_325_b : _GEN_1704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1706 = 9'h146 == r_count_3_io_out ? io_r_326_b : _GEN_1705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1707 = 9'h147 == r_count_3_io_out ? io_r_327_b : _GEN_1706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1708 = 9'h148 == r_count_3_io_out ? io_r_328_b : _GEN_1707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1709 = 9'h149 == r_count_3_io_out ? io_r_329_b : _GEN_1708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1710 = 9'h14a == r_count_3_io_out ? io_r_330_b : _GEN_1709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1711 = 9'h14b == r_count_3_io_out ? io_r_331_b : _GEN_1710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1712 = 9'h14c == r_count_3_io_out ? io_r_332_b : _GEN_1711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1713 = 9'h14d == r_count_3_io_out ? io_r_333_b : _GEN_1712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1714 = 9'h14e == r_count_3_io_out ? io_r_334_b : _GEN_1713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1715 = 9'h14f == r_count_3_io_out ? io_r_335_b : _GEN_1714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1716 = 9'h150 == r_count_3_io_out ? io_r_336_b : _GEN_1715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1717 = 9'h151 == r_count_3_io_out ? io_r_337_b : _GEN_1716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1718 = 9'h152 == r_count_3_io_out ? io_r_338_b : _GEN_1717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1719 = 9'h153 == r_count_3_io_out ? io_r_339_b : _GEN_1718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1720 = 9'h154 == r_count_3_io_out ? io_r_340_b : _GEN_1719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1721 = 9'h155 == r_count_3_io_out ? io_r_341_b : _GEN_1720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1722 = 9'h156 == r_count_3_io_out ? io_r_342_b : _GEN_1721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1723 = 9'h157 == r_count_3_io_out ? io_r_343_b : _GEN_1722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1724 = 9'h158 == r_count_3_io_out ? io_r_344_b : _GEN_1723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1725 = 9'h159 == r_count_3_io_out ? io_r_345_b : _GEN_1724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1726 = 9'h15a == r_count_3_io_out ? io_r_346_b : _GEN_1725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1727 = 9'h15b == r_count_3_io_out ? io_r_347_b : _GEN_1726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1728 = 9'h15c == r_count_3_io_out ? io_r_348_b : _GEN_1727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1729 = 9'h15d == r_count_3_io_out ? io_r_349_b : _GEN_1728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1730 = 9'h15e == r_count_3_io_out ? io_r_350_b : _GEN_1729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1731 = 9'h15f == r_count_3_io_out ? io_r_351_b : _GEN_1730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1732 = 9'h160 == r_count_3_io_out ? io_r_352_b : _GEN_1731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1733 = 9'h161 == r_count_3_io_out ? io_r_353_b : _GEN_1732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1734 = 9'h162 == r_count_3_io_out ? io_r_354_b : _GEN_1733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1735 = 9'h163 == r_count_3_io_out ? io_r_355_b : _GEN_1734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1736 = 9'h164 == r_count_3_io_out ? io_r_356_b : _GEN_1735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1737 = 9'h165 == r_count_3_io_out ? io_r_357_b : _GEN_1736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1738 = 9'h166 == r_count_3_io_out ? io_r_358_b : _GEN_1737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1739 = 9'h167 == r_count_3_io_out ? io_r_359_b : _GEN_1738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1740 = 9'h168 == r_count_3_io_out ? io_r_360_b : _GEN_1739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1741 = 9'h169 == r_count_3_io_out ? io_r_361_b : _GEN_1740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1742 = 9'h16a == r_count_3_io_out ? io_r_362_b : _GEN_1741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1743 = 9'h16b == r_count_3_io_out ? io_r_363_b : _GEN_1742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1744 = 9'h16c == r_count_3_io_out ? io_r_364_b : _GEN_1743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1745 = 9'h16d == r_count_3_io_out ? io_r_365_b : _GEN_1744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1746 = 9'h16e == r_count_3_io_out ? io_r_366_b : _GEN_1745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1747 = 9'h16f == r_count_3_io_out ? io_r_367_b : _GEN_1746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1748 = 9'h170 == r_count_3_io_out ? io_r_368_b : _GEN_1747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1749 = 9'h171 == r_count_3_io_out ? io_r_369_b : _GEN_1748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1750 = 9'h172 == r_count_3_io_out ? io_r_370_b : _GEN_1749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1751 = 9'h173 == r_count_3_io_out ? io_r_371_b : _GEN_1750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1752 = 9'h174 == r_count_3_io_out ? io_r_372_b : _GEN_1751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1753 = 9'h175 == r_count_3_io_out ? io_r_373_b : _GEN_1752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1754 = 9'h176 == r_count_3_io_out ? io_r_374_b : _GEN_1753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1755 = 9'h177 == r_count_3_io_out ? io_r_375_b : _GEN_1754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1756 = 9'h178 == r_count_3_io_out ? io_r_376_b : _GEN_1755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1757 = 9'h179 == r_count_3_io_out ? io_r_377_b : _GEN_1756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1758 = 9'h17a == r_count_3_io_out ? io_r_378_b : _GEN_1757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1759 = 9'h17b == r_count_3_io_out ? io_r_379_b : _GEN_1758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1760 = 9'h17c == r_count_3_io_out ? io_r_380_b : _GEN_1759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1761 = 9'h17d == r_count_3_io_out ? io_r_381_b : _GEN_1760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1762 = 9'h17e == r_count_3_io_out ? io_r_382_b : _GEN_1761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1763 = 9'h17f == r_count_3_io_out ? io_r_383_b : _GEN_1762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1764 = 9'h180 == r_count_3_io_out ? io_r_384_b : _GEN_1763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1765 = 9'h181 == r_count_3_io_out ? io_r_385_b : _GEN_1764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1766 = 9'h182 == r_count_3_io_out ? io_r_386_b : _GEN_1765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1767 = 9'h183 == r_count_3_io_out ? io_r_387_b : _GEN_1766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1768 = 9'h184 == r_count_3_io_out ? io_r_388_b : _GEN_1767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1769 = 9'h185 == r_count_3_io_out ? io_r_389_b : _GEN_1768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1770 = 9'h186 == r_count_3_io_out ? io_r_390_b : _GEN_1769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1771 = 9'h187 == r_count_3_io_out ? io_r_391_b : _GEN_1770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1772 = 9'h188 == r_count_3_io_out ? io_r_392_b : _GEN_1771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1773 = 9'h189 == r_count_3_io_out ? io_r_393_b : _GEN_1772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1774 = 9'h18a == r_count_3_io_out ? io_r_394_b : _GEN_1773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1775 = 9'h18b == r_count_3_io_out ? io_r_395_b : _GEN_1774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1776 = 9'h18c == r_count_3_io_out ? io_r_396_b : _GEN_1775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1777 = 9'h18d == r_count_3_io_out ? io_r_397_b : _GEN_1776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1778 = 9'h18e == r_count_3_io_out ? io_r_398_b : _GEN_1777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1781 = 9'h1 == r_count_4_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1782 = 9'h2 == r_count_4_io_out ? io_r_2_b : _GEN_1781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1783 = 9'h3 == r_count_4_io_out ? io_r_3_b : _GEN_1782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1784 = 9'h4 == r_count_4_io_out ? io_r_4_b : _GEN_1783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1785 = 9'h5 == r_count_4_io_out ? io_r_5_b : _GEN_1784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1786 = 9'h6 == r_count_4_io_out ? io_r_6_b : _GEN_1785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1787 = 9'h7 == r_count_4_io_out ? io_r_7_b : _GEN_1786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1788 = 9'h8 == r_count_4_io_out ? io_r_8_b : _GEN_1787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1789 = 9'h9 == r_count_4_io_out ? io_r_9_b : _GEN_1788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1790 = 9'ha == r_count_4_io_out ? io_r_10_b : _GEN_1789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1791 = 9'hb == r_count_4_io_out ? io_r_11_b : _GEN_1790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1792 = 9'hc == r_count_4_io_out ? io_r_12_b : _GEN_1791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1793 = 9'hd == r_count_4_io_out ? io_r_13_b : _GEN_1792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1794 = 9'he == r_count_4_io_out ? io_r_14_b : _GEN_1793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1795 = 9'hf == r_count_4_io_out ? io_r_15_b : _GEN_1794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1796 = 9'h10 == r_count_4_io_out ? io_r_16_b : _GEN_1795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1797 = 9'h11 == r_count_4_io_out ? io_r_17_b : _GEN_1796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1798 = 9'h12 == r_count_4_io_out ? io_r_18_b : _GEN_1797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1799 = 9'h13 == r_count_4_io_out ? io_r_19_b : _GEN_1798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1800 = 9'h14 == r_count_4_io_out ? io_r_20_b : _GEN_1799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1801 = 9'h15 == r_count_4_io_out ? io_r_21_b : _GEN_1800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1802 = 9'h16 == r_count_4_io_out ? io_r_22_b : _GEN_1801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1803 = 9'h17 == r_count_4_io_out ? io_r_23_b : _GEN_1802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1804 = 9'h18 == r_count_4_io_out ? io_r_24_b : _GEN_1803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1805 = 9'h19 == r_count_4_io_out ? io_r_25_b : _GEN_1804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1806 = 9'h1a == r_count_4_io_out ? io_r_26_b : _GEN_1805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1807 = 9'h1b == r_count_4_io_out ? io_r_27_b : _GEN_1806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1808 = 9'h1c == r_count_4_io_out ? io_r_28_b : _GEN_1807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1809 = 9'h1d == r_count_4_io_out ? io_r_29_b : _GEN_1808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1810 = 9'h1e == r_count_4_io_out ? io_r_30_b : _GEN_1809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1811 = 9'h1f == r_count_4_io_out ? io_r_31_b : _GEN_1810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1812 = 9'h20 == r_count_4_io_out ? io_r_32_b : _GEN_1811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1813 = 9'h21 == r_count_4_io_out ? io_r_33_b : _GEN_1812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1814 = 9'h22 == r_count_4_io_out ? io_r_34_b : _GEN_1813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1815 = 9'h23 == r_count_4_io_out ? io_r_35_b : _GEN_1814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1816 = 9'h24 == r_count_4_io_out ? io_r_36_b : _GEN_1815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1817 = 9'h25 == r_count_4_io_out ? io_r_37_b : _GEN_1816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1818 = 9'h26 == r_count_4_io_out ? io_r_38_b : _GEN_1817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1819 = 9'h27 == r_count_4_io_out ? io_r_39_b : _GEN_1818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1820 = 9'h28 == r_count_4_io_out ? io_r_40_b : _GEN_1819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1821 = 9'h29 == r_count_4_io_out ? io_r_41_b : _GEN_1820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1822 = 9'h2a == r_count_4_io_out ? io_r_42_b : _GEN_1821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1823 = 9'h2b == r_count_4_io_out ? io_r_43_b : _GEN_1822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1824 = 9'h2c == r_count_4_io_out ? io_r_44_b : _GEN_1823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1825 = 9'h2d == r_count_4_io_out ? io_r_45_b : _GEN_1824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1826 = 9'h2e == r_count_4_io_out ? io_r_46_b : _GEN_1825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1827 = 9'h2f == r_count_4_io_out ? io_r_47_b : _GEN_1826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1828 = 9'h30 == r_count_4_io_out ? io_r_48_b : _GEN_1827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1829 = 9'h31 == r_count_4_io_out ? io_r_49_b : _GEN_1828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1830 = 9'h32 == r_count_4_io_out ? io_r_50_b : _GEN_1829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1831 = 9'h33 == r_count_4_io_out ? io_r_51_b : _GEN_1830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1832 = 9'h34 == r_count_4_io_out ? io_r_52_b : _GEN_1831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1833 = 9'h35 == r_count_4_io_out ? io_r_53_b : _GEN_1832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1834 = 9'h36 == r_count_4_io_out ? io_r_54_b : _GEN_1833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1835 = 9'h37 == r_count_4_io_out ? io_r_55_b : _GEN_1834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1836 = 9'h38 == r_count_4_io_out ? io_r_56_b : _GEN_1835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1837 = 9'h39 == r_count_4_io_out ? io_r_57_b : _GEN_1836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1838 = 9'h3a == r_count_4_io_out ? io_r_58_b : _GEN_1837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1839 = 9'h3b == r_count_4_io_out ? io_r_59_b : _GEN_1838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1840 = 9'h3c == r_count_4_io_out ? io_r_60_b : _GEN_1839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1841 = 9'h3d == r_count_4_io_out ? io_r_61_b : _GEN_1840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1842 = 9'h3e == r_count_4_io_out ? io_r_62_b : _GEN_1841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1843 = 9'h3f == r_count_4_io_out ? io_r_63_b : _GEN_1842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1844 = 9'h40 == r_count_4_io_out ? io_r_64_b : _GEN_1843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1845 = 9'h41 == r_count_4_io_out ? io_r_65_b : _GEN_1844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1846 = 9'h42 == r_count_4_io_out ? io_r_66_b : _GEN_1845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1847 = 9'h43 == r_count_4_io_out ? io_r_67_b : _GEN_1846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1848 = 9'h44 == r_count_4_io_out ? io_r_68_b : _GEN_1847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1849 = 9'h45 == r_count_4_io_out ? io_r_69_b : _GEN_1848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1850 = 9'h46 == r_count_4_io_out ? io_r_70_b : _GEN_1849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1851 = 9'h47 == r_count_4_io_out ? io_r_71_b : _GEN_1850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1852 = 9'h48 == r_count_4_io_out ? io_r_72_b : _GEN_1851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1853 = 9'h49 == r_count_4_io_out ? io_r_73_b : _GEN_1852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1854 = 9'h4a == r_count_4_io_out ? io_r_74_b : _GEN_1853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1855 = 9'h4b == r_count_4_io_out ? io_r_75_b : _GEN_1854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1856 = 9'h4c == r_count_4_io_out ? io_r_76_b : _GEN_1855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1857 = 9'h4d == r_count_4_io_out ? io_r_77_b : _GEN_1856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1858 = 9'h4e == r_count_4_io_out ? io_r_78_b : _GEN_1857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1859 = 9'h4f == r_count_4_io_out ? io_r_79_b : _GEN_1858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1860 = 9'h50 == r_count_4_io_out ? io_r_80_b : _GEN_1859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1861 = 9'h51 == r_count_4_io_out ? io_r_81_b : _GEN_1860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1862 = 9'h52 == r_count_4_io_out ? io_r_82_b : _GEN_1861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1863 = 9'h53 == r_count_4_io_out ? io_r_83_b : _GEN_1862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1864 = 9'h54 == r_count_4_io_out ? io_r_84_b : _GEN_1863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1865 = 9'h55 == r_count_4_io_out ? io_r_85_b : _GEN_1864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1866 = 9'h56 == r_count_4_io_out ? io_r_86_b : _GEN_1865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1867 = 9'h57 == r_count_4_io_out ? io_r_87_b : _GEN_1866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1868 = 9'h58 == r_count_4_io_out ? io_r_88_b : _GEN_1867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1869 = 9'h59 == r_count_4_io_out ? io_r_89_b : _GEN_1868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1870 = 9'h5a == r_count_4_io_out ? io_r_90_b : _GEN_1869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1871 = 9'h5b == r_count_4_io_out ? io_r_91_b : _GEN_1870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1872 = 9'h5c == r_count_4_io_out ? io_r_92_b : _GEN_1871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1873 = 9'h5d == r_count_4_io_out ? io_r_93_b : _GEN_1872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1874 = 9'h5e == r_count_4_io_out ? io_r_94_b : _GEN_1873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1875 = 9'h5f == r_count_4_io_out ? io_r_95_b : _GEN_1874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1876 = 9'h60 == r_count_4_io_out ? io_r_96_b : _GEN_1875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1877 = 9'h61 == r_count_4_io_out ? io_r_97_b : _GEN_1876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1878 = 9'h62 == r_count_4_io_out ? io_r_98_b : _GEN_1877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1879 = 9'h63 == r_count_4_io_out ? io_r_99_b : _GEN_1878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1880 = 9'h64 == r_count_4_io_out ? io_r_100_b : _GEN_1879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1881 = 9'h65 == r_count_4_io_out ? io_r_101_b : _GEN_1880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1882 = 9'h66 == r_count_4_io_out ? io_r_102_b : _GEN_1881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1883 = 9'h67 == r_count_4_io_out ? io_r_103_b : _GEN_1882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1884 = 9'h68 == r_count_4_io_out ? io_r_104_b : _GEN_1883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1885 = 9'h69 == r_count_4_io_out ? io_r_105_b : _GEN_1884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1886 = 9'h6a == r_count_4_io_out ? io_r_106_b : _GEN_1885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1887 = 9'h6b == r_count_4_io_out ? io_r_107_b : _GEN_1886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1888 = 9'h6c == r_count_4_io_out ? io_r_108_b : _GEN_1887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1889 = 9'h6d == r_count_4_io_out ? io_r_109_b : _GEN_1888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1890 = 9'h6e == r_count_4_io_out ? io_r_110_b : _GEN_1889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1891 = 9'h6f == r_count_4_io_out ? io_r_111_b : _GEN_1890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1892 = 9'h70 == r_count_4_io_out ? io_r_112_b : _GEN_1891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1893 = 9'h71 == r_count_4_io_out ? io_r_113_b : _GEN_1892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1894 = 9'h72 == r_count_4_io_out ? io_r_114_b : _GEN_1893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1895 = 9'h73 == r_count_4_io_out ? io_r_115_b : _GEN_1894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1896 = 9'h74 == r_count_4_io_out ? io_r_116_b : _GEN_1895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1897 = 9'h75 == r_count_4_io_out ? io_r_117_b : _GEN_1896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1898 = 9'h76 == r_count_4_io_out ? io_r_118_b : _GEN_1897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1899 = 9'h77 == r_count_4_io_out ? io_r_119_b : _GEN_1898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1900 = 9'h78 == r_count_4_io_out ? io_r_120_b : _GEN_1899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1901 = 9'h79 == r_count_4_io_out ? io_r_121_b : _GEN_1900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1902 = 9'h7a == r_count_4_io_out ? io_r_122_b : _GEN_1901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1903 = 9'h7b == r_count_4_io_out ? io_r_123_b : _GEN_1902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1904 = 9'h7c == r_count_4_io_out ? io_r_124_b : _GEN_1903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1905 = 9'h7d == r_count_4_io_out ? io_r_125_b : _GEN_1904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1906 = 9'h7e == r_count_4_io_out ? io_r_126_b : _GEN_1905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1907 = 9'h7f == r_count_4_io_out ? io_r_127_b : _GEN_1906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1908 = 9'h80 == r_count_4_io_out ? io_r_128_b : _GEN_1907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1909 = 9'h81 == r_count_4_io_out ? io_r_129_b : _GEN_1908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1910 = 9'h82 == r_count_4_io_out ? io_r_130_b : _GEN_1909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1911 = 9'h83 == r_count_4_io_out ? io_r_131_b : _GEN_1910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1912 = 9'h84 == r_count_4_io_out ? io_r_132_b : _GEN_1911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1913 = 9'h85 == r_count_4_io_out ? io_r_133_b : _GEN_1912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1914 = 9'h86 == r_count_4_io_out ? io_r_134_b : _GEN_1913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1915 = 9'h87 == r_count_4_io_out ? io_r_135_b : _GEN_1914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1916 = 9'h88 == r_count_4_io_out ? io_r_136_b : _GEN_1915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1917 = 9'h89 == r_count_4_io_out ? io_r_137_b : _GEN_1916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1918 = 9'h8a == r_count_4_io_out ? io_r_138_b : _GEN_1917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1919 = 9'h8b == r_count_4_io_out ? io_r_139_b : _GEN_1918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1920 = 9'h8c == r_count_4_io_out ? io_r_140_b : _GEN_1919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1921 = 9'h8d == r_count_4_io_out ? io_r_141_b : _GEN_1920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1922 = 9'h8e == r_count_4_io_out ? io_r_142_b : _GEN_1921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1923 = 9'h8f == r_count_4_io_out ? io_r_143_b : _GEN_1922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1924 = 9'h90 == r_count_4_io_out ? io_r_144_b : _GEN_1923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1925 = 9'h91 == r_count_4_io_out ? io_r_145_b : _GEN_1924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1926 = 9'h92 == r_count_4_io_out ? io_r_146_b : _GEN_1925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1927 = 9'h93 == r_count_4_io_out ? io_r_147_b : _GEN_1926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1928 = 9'h94 == r_count_4_io_out ? io_r_148_b : _GEN_1927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1929 = 9'h95 == r_count_4_io_out ? io_r_149_b : _GEN_1928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1930 = 9'h96 == r_count_4_io_out ? io_r_150_b : _GEN_1929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1931 = 9'h97 == r_count_4_io_out ? io_r_151_b : _GEN_1930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1932 = 9'h98 == r_count_4_io_out ? io_r_152_b : _GEN_1931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1933 = 9'h99 == r_count_4_io_out ? io_r_153_b : _GEN_1932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1934 = 9'h9a == r_count_4_io_out ? io_r_154_b : _GEN_1933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1935 = 9'h9b == r_count_4_io_out ? io_r_155_b : _GEN_1934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1936 = 9'h9c == r_count_4_io_out ? io_r_156_b : _GEN_1935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1937 = 9'h9d == r_count_4_io_out ? io_r_157_b : _GEN_1936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1938 = 9'h9e == r_count_4_io_out ? io_r_158_b : _GEN_1937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1939 = 9'h9f == r_count_4_io_out ? io_r_159_b : _GEN_1938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1940 = 9'ha0 == r_count_4_io_out ? io_r_160_b : _GEN_1939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1941 = 9'ha1 == r_count_4_io_out ? io_r_161_b : _GEN_1940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1942 = 9'ha2 == r_count_4_io_out ? io_r_162_b : _GEN_1941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1943 = 9'ha3 == r_count_4_io_out ? io_r_163_b : _GEN_1942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1944 = 9'ha4 == r_count_4_io_out ? io_r_164_b : _GEN_1943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1945 = 9'ha5 == r_count_4_io_out ? io_r_165_b : _GEN_1944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1946 = 9'ha6 == r_count_4_io_out ? io_r_166_b : _GEN_1945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1947 = 9'ha7 == r_count_4_io_out ? io_r_167_b : _GEN_1946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1948 = 9'ha8 == r_count_4_io_out ? io_r_168_b : _GEN_1947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1949 = 9'ha9 == r_count_4_io_out ? io_r_169_b : _GEN_1948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1950 = 9'haa == r_count_4_io_out ? io_r_170_b : _GEN_1949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1951 = 9'hab == r_count_4_io_out ? io_r_171_b : _GEN_1950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1952 = 9'hac == r_count_4_io_out ? io_r_172_b : _GEN_1951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1953 = 9'had == r_count_4_io_out ? io_r_173_b : _GEN_1952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1954 = 9'hae == r_count_4_io_out ? io_r_174_b : _GEN_1953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1955 = 9'haf == r_count_4_io_out ? io_r_175_b : _GEN_1954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1956 = 9'hb0 == r_count_4_io_out ? io_r_176_b : _GEN_1955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1957 = 9'hb1 == r_count_4_io_out ? io_r_177_b : _GEN_1956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1958 = 9'hb2 == r_count_4_io_out ? io_r_178_b : _GEN_1957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1959 = 9'hb3 == r_count_4_io_out ? io_r_179_b : _GEN_1958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1960 = 9'hb4 == r_count_4_io_out ? io_r_180_b : _GEN_1959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1961 = 9'hb5 == r_count_4_io_out ? io_r_181_b : _GEN_1960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1962 = 9'hb6 == r_count_4_io_out ? io_r_182_b : _GEN_1961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1963 = 9'hb7 == r_count_4_io_out ? io_r_183_b : _GEN_1962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1964 = 9'hb8 == r_count_4_io_out ? io_r_184_b : _GEN_1963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1965 = 9'hb9 == r_count_4_io_out ? io_r_185_b : _GEN_1964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1966 = 9'hba == r_count_4_io_out ? io_r_186_b : _GEN_1965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1967 = 9'hbb == r_count_4_io_out ? io_r_187_b : _GEN_1966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1968 = 9'hbc == r_count_4_io_out ? io_r_188_b : _GEN_1967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1969 = 9'hbd == r_count_4_io_out ? io_r_189_b : _GEN_1968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1970 = 9'hbe == r_count_4_io_out ? io_r_190_b : _GEN_1969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1971 = 9'hbf == r_count_4_io_out ? io_r_191_b : _GEN_1970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1972 = 9'hc0 == r_count_4_io_out ? io_r_192_b : _GEN_1971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1973 = 9'hc1 == r_count_4_io_out ? io_r_193_b : _GEN_1972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1974 = 9'hc2 == r_count_4_io_out ? io_r_194_b : _GEN_1973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1975 = 9'hc3 == r_count_4_io_out ? io_r_195_b : _GEN_1974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1976 = 9'hc4 == r_count_4_io_out ? io_r_196_b : _GEN_1975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1977 = 9'hc5 == r_count_4_io_out ? io_r_197_b : _GEN_1976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1978 = 9'hc6 == r_count_4_io_out ? io_r_198_b : _GEN_1977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1979 = 9'hc7 == r_count_4_io_out ? io_r_199_b : _GEN_1978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1980 = 9'hc8 == r_count_4_io_out ? io_r_200_b : _GEN_1979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1981 = 9'hc9 == r_count_4_io_out ? io_r_201_b : _GEN_1980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1982 = 9'hca == r_count_4_io_out ? io_r_202_b : _GEN_1981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1983 = 9'hcb == r_count_4_io_out ? io_r_203_b : _GEN_1982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1984 = 9'hcc == r_count_4_io_out ? io_r_204_b : _GEN_1983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1985 = 9'hcd == r_count_4_io_out ? io_r_205_b : _GEN_1984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1986 = 9'hce == r_count_4_io_out ? io_r_206_b : _GEN_1985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1987 = 9'hcf == r_count_4_io_out ? io_r_207_b : _GEN_1986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1988 = 9'hd0 == r_count_4_io_out ? io_r_208_b : _GEN_1987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1989 = 9'hd1 == r_count_4_io_out ? io_r_209_b : _GEN_1988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1990 = 9'hd2 == r_count_4_io_out ? io_r_210_b : _GEN_1989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1991 = 9'hd3 == r_count_4_io_out ? io_r_211_b : _GEN_1990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1992 = 9'hd4 == r_count_4_io_out ? io_r_212_b : _GEN_1991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1993 = 9'hd5 == r_count_4_io_out ? io_r_213_b : _GEN_1992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1994 = 9'hd6 == r_count_4_io_out ? io_r_214_b : _GEN_1993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1995 = 9'hd7 == r_count_4_io_out ? io_r_215_b : _GEN_1994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1996 = 9'hd8 == r_count_4_io_out ? io_r_216_b : _GEN_1995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1997 = 9'hd9 == r_count_4_io_out ? io_r_217_b : _GEN_1996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1998 = 9'hda == r_count_4_io_out ? io_r_218_b : _GEN_1997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1999 = 9'hdb == r_count_4_io_out ? io_r_219_b : _GEN_1998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2000 = 9'hdc == r_count_4_io_out ? io_r_220_b : _GEN_1999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2001 = 9'hdd == r_count_4_io_out ? io_r_221_b : _GEN_2000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2002 = 9'hde == r_count_4_io_out ? io_r_222_b : _GEN_2001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2003 = 9'hdf == r_count_4_io_out ? io_r_223_b : _GEN_2002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2004 = 9'he0 == r_count_4_io_out ? io_r_224_b : _GEN_2003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2005 = 9'he1 == r_count_4_io_out ? io_r_225_b : _GEN_2004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2006 = 9'he2 == r_count_4_io_out ? io_r_226_b : _GEN_2005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2007 = 9'he3 == r_count_4_io_out ? io_r_227_b : _GEN_2006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2008 = 9'he4 == r_count_4_io_out ? io_r_228_b : _GEN_2007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2009 = 9'he5 == r_count_4_io_out ? io_r_229_b : _GEN_2008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2010 = 9'he6 == r_count_4_io_out ? io_r_230_b : _GEN_2009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2011 = 9'he7 == r_count_4_io_out ? io_r_231_b : _GEN_2010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2012 = 9'he8 == r_count_4_io_out ? io_r_232_b : _GEN_2011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2013 = 9'he9 == r_count_4_io_out ? io_r_233_b : _GEN_2012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2014 = 9'hea == r_count_4_io_out ? io_r_234_b : _GEN_2013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2015 = 9'heb == r_count_4_io_out ? io_r_235_b : _GEN_2014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2016 = 9'hec == r_count_4_io_out ? io_r_236_b : _GEN_2015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2017 = 9'hed == r_count_4_io_out ? io_r_237_b : _GEN_2016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2018 = 9'hee == r_count_4_io_out ? io_r_238_b : _GEN_2017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2019 = 9'hef == r_count_4_io_out ? io_r_239_b : _GEN_2018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2020 = 9'hf0 == r_count_4_io_out ? io_r_240_b : _GEN_2019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2021 = 9'hf1 == r_count_4_io_out ? io_r_241_b : _GEN_2020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2022 = 9'hf2 == r_count_4_io_out ? io_r_242_b : _GEN_2021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2023 = 9'hf3 == r_count_4_io_out ? io_r_243_b : _GEN_2022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2024 = 9'hf4 == r_count_4_io_out ? io_r_244_b : _GEN_2023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2025 = 9'hf5 == r_count_4_io_out ? io_r_245_b : _GEN_2024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2026 = 9'hf6 == r_count_4_io_out ? io_r_246_b : _GEN_2025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2027 = 9'hf7 == r_count_4_io_out ? io_r_247_b : _GEN_2026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2028 = 9'hf8 == r_count_4_io_out ? io_r_248_b : _GEN_2027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2029 = 9'hf9 == r_count_4_io_out ? io_r_249_b : _GEN_2028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2030 = 9'hfa == r_count_4_io_out ? io_r_250_b : _GEN_2029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2031 = 9'hfb == r_count_4_io_out ? io_r_251_b : _GEN_2030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2032 = 9'hfc == r_count_4_io_out ? io_r_252_b : _GEN_2031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2033 = 9'hfd == r_count_4_io_out ? io_r_253_b : _GEN_2032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2034 = 9'hfe == r_count_4_io_out ? io_r_254_b : _GEN_2033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2035 = 9'hff == r_count_4_io_out ? io_r_255_b : _GEN_2034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2036 = 9'h100 == r_count_4_io_out ? io_r_256_b : _GEN_2035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2037 = 9'h101 == r_count_4_io_out ? io_r_257_b : _GEN_2036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2038 = 9'h102 == r_count_4_io_out ? io_r_258_b : _GEN_2037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2039 = 9'h103 == r_count_4_io_out ? io_r_259_b : _GEN_2038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2040 = 9'h104 == r_count_4_io_out ? io_r_260_b : _GEN_2039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2041 = 9'h105 == r_count_4_io_out ? io_r_261_b : _GEN_2040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2042 = 9'h106 == r_count_4_io_out ? io_r_262_b : _GEN_2041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2043 = 9'h107 == r_count_4_io_out ? io_r_263_b : _GEN_2042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2044 = 9'h108 == r_count_4_io_out ? io_r_264_b : _GEN_2043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2045 = 9'h109 == r_count_4_io_out ? io_r_265_b : _GEN_2044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2046 = 9'h10a == r_count_4_io_out ? io_r_266_b : _GEN_2045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2047 = 9'h10b == r_count_4_io_out ? io_r_267_b : _GEN_2046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2048 = 9'h10c == r_count_4_io_out ? io_r_268_b : _GEN_2047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2049 = 9'h10d == r_count_4_io_out ? io_r_269_b : _GEN_2048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2050 = 9'h10e == r_count_4_io_out ? io_r_270_b : _GEN_2049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2051 = 9'h10f == r_count_4_io_out ? io_r_271_b : _GEN_2050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2052 = 9'h110 == r_count_4_io_out ? io_r_272_b : _GEN_2051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2053 = 9'h111 == r_count_4_io_out ? io_r_273_b : _GEN_2052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2054 = 9'h112 == r_count_4_io_out ? io_r_274_b : _GEN_2053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2055 = 9'h113 == r_count_4_io_out ? io_r_275_b : _GEN_2054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2056 = 9'h114 == r_count_4_io_out ? io_r_276_b : _GEN_2055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2057 = 9'h115 == r_count_4_io_out ? io_r_277_b : _GEN_2056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2058 = 9'h116 == r_count_4_io_out ? io_r_278_b : _GEN_2057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2059 = 9'h117 == r_count_4_io_out ? io_r_279_b : _GEN_2058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2060 = 9'h118 == r_count_4_io_out ? io_r_280_b : _GEN_2059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2061 = 9'h119 == r_count_4_io_out ? io_r_281_b : _GEN_2060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2062 = 9'h11a == r_count_4_io_out ? io_r_282_b : _GEN_2061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2063 = 9'h11b == r_count_4_io_out ? io_r_283_b : _GEN_2062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2064 = 9'h11c == r_count_4_io_out ? io_r_284_b : _GEN_2063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2065 = 9'h11d == r_count_4_io_out ? io_r_285_b : _GEN_2064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2066 = 9'h11e == r_count_4_io_out ? io_r_286_b : _GEN_2065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2067 = 9'h11f == r_count_4_io_out ? io_r_287_b : _GEN_2066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2068 = 9'h120 == r_count_4_io_out ? io_r_288_b : _GEN_2067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2069 = 9'h121 == r_count_4_io_out ? io_r_289_b : _GEN_2068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2070 = 9'h122 == r_count_4_io_out ? io_r_290_b : _GEN_2069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2071 = 9'h123 == r_count_4_io_out ? io_r_291_b : _GEN_2070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2072 = 9'h124 == r_count_4_io_out ? io_r_292_b : _GEN_2071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2073 = 9'h125 == r_count_4_io_out ? io_r_293_b : _GEN_2072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2074 = 9'h126 == r_count_4_io_out ? io_r_294_b : _GEN_2073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2075 = 9'h127 == r_count_4_io_out ? io_r_295_b : _GEN_2074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2076 = 9'h128 == r_count_4_io_out ? io_r_296_b : _GEN_2075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2077 = 9'h129 == r_count_4_io_out ? io_r_297_b : _GEN_2076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2078 = 9'h12a == r_count_4_io_out ? io_r_298_b : _GEN_2077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2079 = 9'h12b == r_count_4_io_out ? io_r_299_b : _GEN_2078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2080 = 9'h12c == r_count_4_io_out ? io_r_300_b : _GEN_2079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2081 = 9'h12d == r_count_4_io_out ? io_r_301_b : _GEN_2080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2082 = 9'h12e == r_count_4_io_out ? io_r_302_b : _GEN_2081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2083 = 9'h12f == r_count_4_io_out ? io_r_303_b : _GEN_2082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2084 = 9'h130 == r_count_4_io_out ? io_r_304_b : _GEN_2083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2085 = 9'h131 == r_count_4_io_out ? io_r_305_b : _GEN_2084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2086 = 9'h132 == r_count_4_io_out ? io_r_306_b : _GEN_2085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2087 = 9'h133 == r_count_4_io_out ? io_r_307_b : _GEN_2086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2088 = 9'h134 == r_count_4_io_out ? io_r_308_b : _GEN_2087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2089 = 9'h135 == r_count_4_io_out ? io_r_309_b : _GEN_2088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2090 = 9'h136 == r_count_4_io_out ? io_r_310_b : _GEN_2089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2091 = 9'h137 == r_count_4_io_out ? io_r_311_b : _GEN_2090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2092 = 9'h138 == r_count_4_io_out ? io_r_312_b : _GEN_2091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2093 = 9'h139 == r_count_4_io_out ? io_r_313_b : _GEN_2092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2094 = 9'h13a == r_count_4_io_out ? io_r_314_b : _GEN_2093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2095 = 9'h13b == r_count_4_io_out ? io_r_315_b : _GEN_2094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2096 = 9'h13c == r_count_4_io_out ? io_r_316_b : _GEN_2095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2097 = 9'h13d == r_count_4_io_out ? io_r_317_b : _GEN_2096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2098 = 9'h13e == r_count_4_io_out ? io_r_318_b : _GEN_2097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2099 = 9'h13f == r_count_4_io_out ? io_r_319_b : _GEN_2098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2100 = 9'h140 == r_count_4_io_out ? io_r_320_b : _GEN_2099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2101 = 9'h141 == r_count_4_io_out ? io_r_321_b : _GEN_2100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2102 = 9'h142 == r_count_4_io_out ? io_r_322_b : _GEN_2101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2103 = 9'h143 == r_count_4_io_out ? io_r_323_b : _GEN_2102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2104 = 9'h144 == r_count_4_io_out ? io_r_324_b : _GEN_2103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2105 = 9'h145 == r_count_4_io_out ? io_r_325_b : _GEN_2104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2106 = 9'h146 == r_count_4_io_out ? io_r_326_b : _GEN_2105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2107 = 9'h147 == r_count_4_io_out ? io_r_327_b : _GEN_2106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2108 = 9'h148 == r_count_4_io_out ? io_r_328_b : _GEN_2107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2109 = 9'h149 == r_count_4_io_out ? io_r_329_b : _GEN_2108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2110 = 9'h14a == r_count_4_io_out ? io_r_330_b : _GEN_2109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2111 = 9'h14b == r_count_4_io_out ? io_r_331_b : _GEN_2110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2112 = 9'h14c == r_count_4_io_out ? io_r_332_b : _GEN_2111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2113 = 9'h14d == r_count_4_io_out ? io_r_333_b : _GEN_2112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2114 = 9'h14e == r_count_4_io_out ? io_r_334_b : _GEN_2113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2115 = 9'h14f == r_count_4_io_out ? io_r_335_b : _GEN_2114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2116 = 9'h150 == r_count_4_io_out ? io_r_336_b : _GEN_2115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2117 = 9'h151 == r_count_4_io_out ? io_r_337_b : _GEN_2116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2118 = 9'h152 == r_count_4_io_out ? io_r_338_b : _GEN_2117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2119 = 9'h153 == r_count_4_io_out ? io_r_339_b : _GEN_2118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2120 = 9'h154 == r_count_4_io_out ? io_r_340_b : _GEN_2119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2121 = 9'h155 == r_count_4_io_out ? io_r_341_b : _GEN_2120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2122 = 9'h156 == r_count_4_io_out ? io_r_342_b : _GEN_2121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2123 = 9'h157 == r_count_4_io_out ? io_r_343_b : _GEN_2122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2124 = 9'h158 == r_count_4_io_out ? io_r_344_b : _GEN_2123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2125 = 9'h159 == r_count_4_io_out ? io_r_345_b : _GEN_2124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2126 = 9'h15a == r_count_4_io_out ? io_r_346_b : _GEN_2125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2127 = 9'h15b == r_count_4_io_out ? io_r_347_b : _GEN_2126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2128 = 9'h15c == r_count_4_io_out ? io_r_348_b : _GEN_2127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2129 = 9'h15d == r_count_4_io_out ? io_r_349_b : _GEN_2128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2130 = 9'h15e == r_count_4_io_out ? io_r_350_b : _GEN_2129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2131 = 9'h15f == r_count_4_io_out ? io_r_351_b : _GEN_2130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2132 = 9'h160 == r_count_4_io_out ? io_r_352_b : _GEN_2131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2133 = 9'h161 == r_count_4_io_out ? io_r_353_b : _GEN_2132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2134 = 9'h162 == r_count_4_io_out ? io_r_354_b : _GEN_2133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2135 = 9'h163 == r_count_4_io_out ? io_r_355_b : _GEN_2134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2136 = 9'h164 == r_count_4_io_out ? io_r_356_b : _GEN_2135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2137 = 9'h165 == r_count_4_io_out ? io_r_357_b : _GEN_2136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2138 = 9'h166 == r_count_4_io_out ? io_r_358_b : _GEN_2137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2139 = 9'h167 == r_count_4_io_out ? io_r_359_b : _GEN_2138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2140 = 9'h168 == r_count_4_io_out ? io_r_360_b : _GEN_2139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2141 = 9'h169 == r_count_4_io_out ? io_r_361_b : _GEN_2140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2142 = 9'h16a == r_count_4_io_out ? io_r_362_b : _GEN_2141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2143 = 9'h16b == r_count_4_io_out ? io_r_363_b : _GEN_2142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2144 = 9'h16c == r_count_4_io_out ? io_r_364_b : _GEN_2143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2145 = 9'h16d == r_count_4_io_out ? io_r_365_b : _GEN_2144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2146 = 9'h16e == r_count_4_io_out ? io_r_366_b : _GEN_2145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2147 = 9'h16f == r_count_4_io_out ? io_r_367_b : _GEN_2146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2148 = 9'h170 == r_count_4_io_out ? io_r_368_b : _GEN_2147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2149 = 9'h171 == r_count_4_io_out ? io_r_369_b : _GEN_2148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2150 = 9'h172 == r_count_4_io_out ? io_r_370_b : _GEN_2149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2151 = 9'h173 == r_count_4_io_out ? io_r_371_b : _GEN_2150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2152 = 9'h174 == r_count_4_io_out ? io_r_372_b : _GEN_2151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2153 = 9'h175 == r_count_4_io_out ? io_r_373_b : _GEN_2152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2154 = 9'h176 == r_count_4_io_out ? io_r_374_b : _GEN_2153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2155 = 9'h177 == r_count_4_io_out ? io_r_375_b : _GEN_2154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2156 = 9'h178 == r_count_4_io_out ? io_r_376_b : _GEN_2155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2157 = 9'h179 == r_count_4_io_out ? io_r_377_b : _GEN_2156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2158 = 9'h17a == r_count_4_io_out ? io_r_378_b : _GEN_2157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2159 = 9'h17b == r_count_4_io_out ? io_r_379_b : _GEN_2158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2160 = 9'h17c == r_count_4_io_out ? io_r_380_b : _GEN_2159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2161 = 9'h17d == r_count_4_io_out ? io_r_381_b : _GEN_2160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2162 = 9'h17e == r_count_4_io_out ? io_r_382_b : _GEN_2161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2163 = 9'h17f == r_count_4_io_out ? io_r_383_b : _GEN_2162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2164 = 9'h180 == r_count_4_io_out ? io_r_384_b : _GEN_2163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2165 = 9'h181 == r_count_4_io_out ? io_r_385_b : _GEN_2164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2166 = 9'h182 == r_count_4_io_out ? io_r_386_b : _GEN_2165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2167 = 9'h183 == r_count_4_io_out ? io_r_387_b : _GEN_2166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2168 = 9'h184 == r_count_4_io_out ? io_r_388_b : _GEN_2167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2169 = 9'h185 == r_count_4_io_out ? io_r_389_b : _GEN_2168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2170 = 9'h186 == r_count_4_io_out ? io_r_390_b : _GEN_2169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2171 = 9'h187 == r_count_4_io_out ? io_r_391_b : _GEN_2170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2172 = 9'h188 == r_count_4_io_out ? io_r_392_b : _GEN_2171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2173 = 9'h189 == r_count_4_io_out ? io_r_393_b : _GEN_2172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2174 = 9'h18a == r_count_4_io_out ? io_r_394_b : _GEN_2173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2175 = 9'h18b == r_count_4_io_out ? io_r_395_b : _GEN_2174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2176 = 9'h18c == r_count_4_io_out ? io_r_396_b : _GEN_2175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2177 = 9'h18d == r_count_4_io_out ? io_r_397_b : _GEN_2176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2178 = 9'h18e == r_count_4_io_out ? io_r_398_b : _GEN_2177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2181 = 9'h1 == r_count_5_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2182 = 9'h2 == r_count_5_io_out ? io_r_2_b : _GEN_2181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2183 = 9'h3 == r_count_5_io_out ? io_r_3_b : _GEN_2182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2184 = 9'h4 == r_count_5_io_out ? io_r_4_b : _GEN_2183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2185 = 9'h5 == r_count_5_io_out ? io_r_5_b : _GEN_2184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2186 = 9'h6 == r_count_5_io_out ? io_r_6_b : _GEN_2185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2187 = 9'h7 == r_count_5_io_out ? io_r_7_b : _GEN_2186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2188 = 9'h8 == r_count_5_io_out ? io_r_8_b : _GEN_2187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2189 = 9'h9 == r_count_5_io_out ? io_r_9_b : _GEN_2188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2190 = 9'ha == r_count_5_io_out ? io_r_10_b : _GEN_2189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2191 = 9'hb == r_count_5_io_out ? io_r_11_b : _GEN_2190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2192 = 9'hc == r_count_5_io_out ? io_r_12_b : _GEN_2191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2193 = 9'hd == r_count_5_io_out ? io_r_13_b : _GEN_2192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2194 = 9'he == r_count_5_io_out ? io_r_14_b : _GEN_2193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2195 = 9'hf == r_count_5_io_out ? io_r_15_b : _GEN_2194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2196 = 9'h10 == r_count_5_io_out ? io_r_16_b : _GEN_2195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2197 = 9'h11 == r_count_5_io_out ? io_r_17_b : _GEN_2196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2198 = 9'h12 == r_count_5_io_out ? io_r_18_b : _GEN_2197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2199 = 9'h13 == r_count_5_io_out ? io_r_19_b : _GEN_2198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2200 = 9'h14 == r_count_5_io_out ? io_r_20_b : _GEN_2199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2201 = 9'h15 == r_count_5_io_out ? io_r_21_b : _GEN_2200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2202 = 9'h16 == r_count_5_io_out ? io_r_22_b : _GEN_2201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2203 = 9'h17 == r_count_5_io_out ? io_r_23_b : _GEN_2202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2204 = 9'h18 == r_count_5_io_out ? io_r_24_b : _GEN_2203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2205 = 9'h19 == r_count_5_io_out ? io_r_25_b : _GEN_2204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2206 = 9'h1a == r_count_5_io_out ? io_r_26_b : _GEN_2205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2207 = 9'h1b == r_count_5_io_out ? io_r_27_b : _GEN_2206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2208 = 9'h1c == r_count_5_io_out ? io_r_28_b : _GEN_2207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2209 = 9'h1d == r_count_5_io_out ? io_r_29_b : _GEN_2208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2210 = 9'h1e == r_count_5_io_out ? io_r_30_b : _GEN_2209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2211 = 9'h1f == r_count_5_io_out ? io_r_31_b : _GEN_2210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2212 = 9'h20 == r_count_5_io_out ? io_r_32_b : _GEN_2211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2213 = 9'h21 == r_count_5_io_out ? io_r_33_b : _GEN_2212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2214 = 9'h22 == r_count_5_io_out ? io_r_34_b : _GEN_2213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2215 = 9'h23 == r_count_5_io_out ? io_r_35_b : _GEN_2214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2216 = 9'h24 == r_count_5_io_out ? io_r_36_b : _GEN_2215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2217 = 9'h25 == r_count_5_io_out ? io_r_37_b : _GEN_2216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2218 = 9'h26 == r_count_5_io_out ? io_r_38_b : _GEN_2217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2219 = 9'h27 == r_count_5_io_out ? io_r_39_b : _GEN_2218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2220 = 9'h28 == r_count_5_io_out ? io_r_40_b : _GEN_2219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2221 = 9'h29 == r_count_5_io_out ? io_r_41_b : _GEN_2220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2222 = 9'h2a == r_count_5_io_out ? io_r_42_b : _GEN_2221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2223 = 9'h2b == r_count_5_io_out ? io_r_43_b : _GEN_2222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2224 = 9'h2c == r_count_5_io_out ? io_r_44_b : _GEN_2223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2225 = 9'h2d == r_count_5_io_out ? io_r_45_b : _GEN_2224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2226 = 9'h2e == r_count_5_io_out ? io_r_46_b : _GEN_2225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2227 = 9'h2f == r_count_5_io_out ? io_r_47_b : _GEN_2226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2228 = 9'h30 == r_count_5_io_out ? io_r_48_b : _GEN_2227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2229 = 9'h31 == r_count_5_io_out ? io_r_49_b : _GEN_2228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2230 = 9'h32 == r_count_5_io_out ? io_r_50_b : _GEN_2229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2231 = 9'h33 == r_count_5_io_out ? io_r_51_b : _GEN_2230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2232 = 9'h34 == r_count_5_io_out ? io_r_52_b : _GEN_2231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2233 = 9'h35 == r_count_5_io_out ? io_r_53_b : _GEN_2232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2234 = 9'h36 == r_count_5_io_out ? io_r_54_b : _GEN_2233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2235 = 9'h37 == r_count_5_io_out ? io_r_55_b : _GEN_2234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2236 = 9'h38 == r_count_5_io_out ? io_r_56_b : _GEN_2235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2237 = 9'h39 == r_count_5_io_out ? io_r_57_b : _GEN_2236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2238 = 9'h3a == r_count_5_io_out ? io_r_58_b : _GEN_2237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2239 = 9'h3b == r_count_5_io_out ? io_r_59_b : _GEN_2238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2240 = 9'h3c == r_count_5_io_out ? io_r_60_b : _GEN_2239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2241 = 9'h3d == r_count_5_io_out ? io_r_61_b : _GEN_2240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2242 = 9'h3e == r_count_5_io_out ? io_r_62_b : _GEN_2241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2243 = 9'h3f == r_count_5_io_out ? io_r_63_b : _GEN_2242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2244 = 9'h40 == r_count_5_io_out ? io_r_64_b : _GEN_2243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2245 = 9'h41 == r_count_5_io_out ? io_r_65_b : _GEN_2244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2246 = 9'h42 == r_count_5_io_out ? io_r_66_b : _GEN_2245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2247 = 9'h43 == r_count_5_io_out ? io_r_67_b : _GEN_2246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2248 = 9'h44 == r_count_5_io_out ? io_r_68_b : _GEN_2247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2249 = 9'h45 == r_count_5_io_out ? io_r_69_b : _GEN_2248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2250 = 9'h46 == r_count_5_io_out ? io_r_70_b : _GEN_2249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2251 = 9'h47 == r_count_5_io_out ? io_r_71_b : _GEN_2250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2252 = 9'h48 == r_count_5_io_out ? io_r_72_b : _GEN_2251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2253 = 9'h49 == r_count_5_io_out ? io_r_73_b : _GEN_2252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2254 = 9'h4a == r_count_5_io_out ? io_r_74_b : _GEN_2253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2255 = 9'h4b == r_count_5_io_out ? io_r_75_b : _GEN_2254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2256 = 9'h4c == r_count_5_io_out ? io_r_76_b : _GEN_2255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2257 = 9'h4d == r_count_5_io_out ? io_r_77_b : _GEN_2256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2258 = 9'h4e == r_count_5_io_out ? io_r_78_b : _GEN_2257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2259 = 9'h4f == r_count_5_io_out ? io_r_79_b : _GEN_2258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2260 = 9'h50 == r_count_5_io_out ? io_r_80_b : _GEN_2259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2261 = 9'h51 == r_count_5_io_out ? io_r_81_b : _GEN_2260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2262 = 9'h52 == r_count_5_io_out ? io_r_82_b : _GEN_2261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2263 = 9'h53 == r_count_5_io_out ? io_r_83_b : _GEN_2262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2264 = 9'h54 == r_count_5_io_out ? io_r_84_b : _GEN_2263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2265 = 9'h55 == r_count_5_io_out ? io_r_85_b : _GEN_2264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2266 = 9'h56 == r_count_5_io_out ? io_r_86_b : _GEN_2265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2267 = 9'h57 == r_count_5_io_out ? io_r_87_b : _GEN_2266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2268 = 9'h58 == r_count_5_io_out ? io_r_88_b : _GEN_2267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2269 = 9'h59 == r_count_5_io_out ? io_r_89_b : _GEN_2268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2270 = 9'h5a == r_count_5_io_out ? io_r_90_b : _GEN_2269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2271 = 9'h5b == r_count_5_io_out ? io_r_91_b : _GEN_2270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2272 = 9'h5c == r_count_5_io_out ? io_r_92_b : _GEN_2271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2273 = 9'h5d == r_count_5_io_out ? io_r_93_b : _GEN_2272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2274 = 9'h5e == r_count_5_io_out ? io_r_94_b : _GEN_2273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2275 = 9'h5f == r_count_5_io_out ? io_r_95_b : _GEN_2274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2276 = 9'h60 == r_count_5_io_out ? io_r_96_b : _GEN_2275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2277 = 9'h61 == r_count_5_io_out ? io_r_97_b : _GEN_2276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2278 = 9'h62 == r_count_5_io_out ? io_r_98_b : _GEN_2277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2279 = 9'h63 == r_count_5_io_out ? io_r_99_b : _GEN_2278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2280 = 9'h64 == r_count_5_io_out ? io_r_100_b : _GEN_2279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2281 = 9'h65 == r_count_5_io_out ? io_r_101_b : _GEN_2280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2282 = 9'h66 == r_count_5_io_out ? io_r_102_b : _GEN_2281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2283 = 9'h67 == r_count_5_io_out ? io_r_103_b : _GEN_2282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2284 = 9'h68 == r_count_5_io_out ? io_r_104_b : _GEN_2283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2285 = 9'h69 == r_count_5_io_out ? io_r_105_b : _GEN_2284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2286 = 9'h6a == r_count_5_io_out ? io_r_106_b : _GEN_2285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2287 = 9'h6b == r_count_5_io_out ? io_r_107_b : _GEN_2286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2288 = 9'h6c == r_count_5_io_out ? io_r_108_b : _GEN_2287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2289 = 9'h6d == r_count_5_io_out ? io_r_109_b : _GEN_2288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2290 = 9'h6e == r_count_5_io_out ? io_r_110_b : _GEN_2289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2291 = 9'h6f == r_count_5_io_out ? io_r_111_b : _GEN_2290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2292 = 9'h70 == r_count_5_io_out ? io_r_112_b : _GEN_2291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2293 = 9'h71 == r_count_5_io_out ? io_r_113_b : _GEN_2292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2294 = 9'h72 == r_count_5_io_out ? io_r_114_b : _GEN_2293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2295 = 9'h73 == r_count_5_io_out ? io_r_115_b : _GEN_2294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2296 = 9'h74 == r_count_5_io_out ? io_r_116_b : _GEN_2295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2297 = 9'h75 == r_count_5_io_out ? io_r_117_b : _GEN_2296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2298 = 9'h76 == r_count_5_io_out ? io_r_118_b : _GEN_2297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2299 = 9'h77 == r_count_5_io_out ? io_r_119_b : _GEN_2298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2300 = 9'h78 == r_count_5_io_out ? io_r_120_b : _GEN_2299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2301 = 9'h79 == r_count_5_io_out ? io_r_121_b : _GEN_2300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2302 = 9'h7a == r_count_5_io_out ? io_r_122_b : _GEN_2301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2303 = 9'h7b == r_count_5_io_out ? io_r_123_b : _GEN_2302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2304 = 9'h7c == r_count_5_io_out ? io_r_124_b : _GEN_2303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2305 = 9'h7d == r_count_5_io_out ? io_r_125_b : _GEN_2304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2306 = 9'h7e == r_count_5_io_out ? io_r_126_b : _GEN_2305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2307 = 9'h7f == r_count_5_io_out ? io_r_127_b : _GEN_2306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2308 = 9'h80 == r_count_5_io_out ? io_r_128_b : _GEN_2307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2309 = 9'h81 == r_count_5_io_out ? io_r_129_b : _GEN_2308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2310 = 9'h82 == r_count_5_io_out ? io_r_130_b : _GEN_2309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2311 = 9'h83 == r_count_5_io_out ? io_r_131_b : _GEN_2310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2312 = 9'h84 == r_count_5_io_out ? io_r_132_b : _GEN_2311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2313 = 9'h85 == r_count_5_io_out ? io_r_133_b : _GEN_2312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2314 = 9'h86 == r_count_5_io_out ? io_r_134_b : _GEN_2313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2315 = 9'h87 == r_count_5_io_out ? io_r_135_b : _GEN_2314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2316 = 9'h88 == r_count_5_io_out ? io_r_136_b : _GEN_2315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2317 = 9'h89 == r_count_5_io_out ? io_r_137_b : _GEN_2316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2318 = 9'h8a == r_count_5_io_out ? io_r_138_b : _GEN_2317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2319 = 9'h8b == r_count_5_io_out ? io_r_139_b : _GEN_2318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2320 = 9'h8c == r_count_5_io_out ? io_r_140_b : _GEN_2319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2321 = 9'h8d == r_count_5_io_out ? io_r_141_b : _GEN_2320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2322 = 9'h8e == r_count_5_io_out ? io_r_142_b : _GEN_2321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2323 = 9'h8f == r_count_5_io_out ? io_r_143_b : _GEN_2322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2324 = 9'h90 == r_count_5_io_out ? io_r_144_b : _GEN_2323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2325 = 9'h91 == r_count_5_io_out ? io_r_145_b : _GEN_2324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2326 = 9'h92 == r_count_5_io_out ? io_r_146_b : _GEN_2325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2327 = 9'h93 == r_count_5_io_out ? io_r_147_b : _GEN_2326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2328 = 9'h94 == r_count_5_io_out ? io_r_148_b : _GEN_2327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2329 = 9'h95 == r_count_5_io_out ? io_r_149_b : _GEN_2328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2330 = 9'h96 == r_count_5_io_out ? io_r_150_b : _GEN_2329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2331 = 9'h97 == r_count_5_io_out ? io_r_151_b : _GEN_2330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2332 = 9'h98 == r_count_5_io_out ? io_r_152_b : _GEN_2331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2333 = 9'h99 == r_count_5_io_out ? io_r_153_b : _GEN_2332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2334 = 9'h9a == r_count_5_io_out ? io_r_154_b : _GEN_2333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2335 = 9'h9b == r_count_5_io_out ? io_r_155_b : _GEN_2334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2336 = 9'h9c == r_count_5_io_out ? io_r_156_b : _GEN_2335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2337 = 9'h9d == r_count_5_io_out ? io_r_157_b : _GEN_2336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2338 = 9'h9e == r_count_5_io_out ? io_r_158_b : _GEN_2337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2339 = 9'h9f == r_count_5_io_out ? io_r_159_b : _GEN_2338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2340 = 9'ha0 == r_count_5_io_out ? io_r_160_b : _GEN_2339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2341 = 9'ha1 == r_count_5_io_out ? io_r_161_b : _GEN_2340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2342 = 9'ha2 == r_count_5_io_out ? io_r_162_b : _GEN_2341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2343 = 9'ha3 == r_count_5_io_out ? io_r_163_b : _GEN_2342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2344 = 9'ha4 == r_count_5_io_out ? io_r_164_b : _GEN_2343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2345 = 9'ha5 == r_count_5_io_out ? io_r_165_b : _GEN_2344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2346 = 9'ha6 == r_count_5_io_out ? io_r_166_b : _GEN_2345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2347 = 9'ha7 == r_count_5_io_out ? io_r_167_b : _GEN_2346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2348 = 9'ha8 == r_count_5_io_out ? io_r_168_b : _GEN_2347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2349 = 9'ha9 == r_count_5_io_out ? io_r_169_b : _GEN_2348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2350 = 9'haa == r_count_5_io_out ? io_r_170_b : _GEN_2349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2351 = 9'hab == r_count_5_io_out ? io_r_171_b : _GEN_2350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2352 = 9'hac == r_count_5_io_out ? io_r_172_b : _GEN_2351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2353 = 9'had == r_count_5_io_out ? io_r_173_b : _GEN_2352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2354 = 9'hae == r_count_5_io_out ? io_r_174_b : _GEN_2353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2355 = 9'haf == r_count_5_io_out ? io_r_175_b : _GEN_2354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2356 = 9'hb0 == r_count_5_io_out ? io_r_176_b : _GEN_2355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2357 = 9'hb1 == r_count_5_io_out ? io_r_177_b : _GEN_2356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2358 = 9'hb2 == r_count_5_io_out ? io_r_178_b : _GEN_2357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2359 = 9'hb3 == r_count_5_io_out ? io_r_179_b : _GEN_2358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2360 = 9'hb4 == r_count_5_io_out ? io_r_180_b : _GEN_2359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2361 = 9'hb5 == r_count_5_io_out ? io_r_181_b : _GEN_2360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2362 = 9'hb6 == r_count_5_io_out ? io_r_182_b : _GEN_2361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2363 = 9'hb7 == r_count_5_io_out ? io_r_183_b : _GEN_2362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2364 = 9'hb8 == r_count_5_io_out ? io_r_184_b : _GEN_2363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2365 = 9'hb9 == r_count_5_io_out ? io_r_185_b : _GEN_2364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2366 = 9'hba == r_count_5_io_out ? io_r_186_b : _GEN_2365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2367 = 9'hbb == r_count_5_io_out ? io_r_187_b : _GEN_2366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2368 = 9'hbc == r_count_5_io_out ? io_r_188_b : _GEN_2367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2369 = 9'hbd == r_count_5_io_out ? io_r_189_b : _GEN_2368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2370 = 9'hbe == r_count_5_io_out ? io_r_190_b : _GEN_2369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2371 = 9'hbf == r_count_5_io_out ? io_r_191_b : _GEN_2370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2372 = 9'hc0 == r_count_5_io_out ? io_r_192_b : _GEN_2371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2373 = 9'hc1 == r_count_5_io_out ? io_r_193_b : _GEN_2372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2374 = 9'hc2 == r_count_5_io_out ? io_r_194_b : _GEN_2373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2375 = 9'hc3 == r_count_5_io_out ? io_r_195_b : _GEN_2374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2376 = 9'hc4 == r_count_5_io_out ? io_r_196_b : _GEN_2375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2377 = 9'hc5 == r_count_5_io_out ? io_r_197_b : _GEN_2376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2378 = 9'hc6 == r_count_5_io_out ? io_r_198_b : _GEN_2377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2379 = 9'hc7 == r_count_5_io_out ? io_r_199_b : _GEN_2378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2380 = 9'hc8 == r_count_5_io_out ? io_r_200_b : _GEN_2379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2381 = 9'hc9 == r_count_5_io_out ? io_r_201_b : _GEN_2380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2382 = 9'hca == r_count_5_io_out ? io_r_202_b : _GEN_2381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2383 = 9'hcb == r_count_5_io_out ? io_r_203_b : _GEN_2382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2384 = 9'hcc == r_count_5_io_out ? io_r_204_b : _GEN_2383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2385 = 9'hcd == r_count_5_io_out ? io_r_205_b : _GEN_2384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2386 = 9'hce == r_count_5_io_out ? io_r_206_b : _GEN_2385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2387 = 9'hcf == r_count_5_io_out ? io_r_207_b : _GEN_2386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2388 = 9'hd0 == r_count_5_io_out ? io_r_208_b : _GEN_2387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2389 = 9'hd1 == r_count_5_io_out ? io_r_209_b : _GEN_2388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2390 = 9'hd2 == r_count_5_io_out ? io_r_210_b : _GEN_2389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2391 = 9'hd3 == r_count_5_io_out ? io_r_211_b : _GEN_2390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2392 = 9'hd4 == r_count_5_io_out ? io_r_212_b : _GEN_2391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2393 = 9'hd5 == r_count_5_io_out ? io_r_213_b : _GEN_2392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2394 = 9'hd6 == r_count_5_io_out ? io_r_214_b : _GEN_2393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2395 = 9'hd7 == r_count_5_io_out ? io_r_215_b : _GEN_2394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2396 = 9'hd8 == r_count_5_io_out ? io_r_216_b : _GEN_2395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2397 = 9'hd9 == r_count_5_io_out ? io_r_217_b : _GEN_2396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2398 = 9'hda == r_count_5_io_out ? io_r_218_b : _GEN_2397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2399 = 9'hdb == r_count_5_io_out ? io_r_219_b : _GEN_2398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2400 = 9'hdc == r_count_5_io_out ? io_r_220_b : _GEN_2399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2401 = 9'hdd == r_count_5_io_out ? io_r_221_b : _GEN_2400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2402 = 9'hde == r_count_5_io_out ? io_r_222_b : _GEN_2401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2403 = 9'hdf == r_count_5_io_out ? io_r_223_b : _GEN_2402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2404 = 9'he0 == r_count_5_io_out ? io_r_224_b : _GEN_2403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2405 = 9'he1 == r_count_5_io_out ? io_r_225_b : _GEN_2404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2406 = 9'he2 == r_count_5_io_out ? io_r_226_b : _GEN_2405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2407 = 9'he3 == r_count_5_io_out ? io_r_227_b : _GEN_2406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2408 = 9'he4 == r_count_5_io_out ? io_r_228_b : _GEN_2407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2409 = 9'he5 == r_count_5_io_out ? io_r_229_b : _GEN_2408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2410 = 9'he6 == r_count_5_io_out ? io_r_230_b : _GEN_2409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2411 = 9'he7 == r_count_5_io_out ? io_r_231_b : _GEN_2410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2412 = 9'he8 == r_count_5_io_out ? io_r_232_b : _GEN_2411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2413 = 9'he9 == r_count_5_io_out ? io_r_233_b : _GEN_2412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2414 = 9'hea == r_count_5_io_out ? io_r_234_b : _GEN_2413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2415 = 9'heb == r_count_5_io_out ? io_r_235_b : _GEN_2414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2416 = 9'hec == r_count_5_io_out ? io_r_236_b : _GEN_2415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2417 = 9'hed == r_count_5_io_out ? io_r_237_b : _GEN_2416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2418 = 9'hee == r_count_5_io_out ? io_r_238_b : _GEN_2417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2419 = 9'hef == r_count_5_io_out ? io_r_239_b : _GEN_2418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2420 = 9'hf0 == r_count_5_io_out ? io_r_240_b : _GEN_2419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2421 = 9'hf1 == r_count_5_io_out ? io_r_241_b : _GEN_2420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2422 = 9'hf2 == r_count_5_io_out ? io_r_242_b : _GEN_2421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2423 = 9'hf3 == r_count_5_io_out ? io_r_243_b : _GEN_2422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2424 = 9'hf4 == r_count_5_io_out ? io_r_244_b : _GEN_2423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2425 = 9'hf5 == r_count_5_io_out ? io_r_245_b : _GEN_2424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2426 = 9'hf6 == r_count_5_io_out ? io_r_246_b : _GEN_2425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2427 = 9'hf7 == r_count_5_io_out ? io_r_247_b : _GEN_2426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2428 = 9'hf8 == r_count_5_io_out ? io_r_248_b : _GEN_2427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2429 = 9'hf9 == r_count_5_io_out ? io_r_249_b : _GEN_2428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2430 = 9'hfa == r_count_5_io_out ? io_r_250_b : _GEN_2429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2431 = 9'hfb == r_count_5_io_out ? io_r_251_b : _GEN_2430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2432 = 9'hfc == r_count_5_io_out ? io_r_252_b : _GEN_2431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2433 = 9'hfd == r_count_5_io_out ? io_r_253_b : _GEN_2432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2434 = 9'hfe == r_count_5_io_out ? io_r_254_b : _GEN_2433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2435 = 9'hff == r_count_5_io_out ? io_r_255_b : _GEN_2434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2436 = 9'h100 == r_count_5_io_out ? io_r_256_b : _GEN_2435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2437 = 9'h101 == r_count_5_io_out ? io_r_257_b : _GEN_2436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2438 = 9'h102 == r_count_5_io_out ? io_r_258_b : _GEN_2437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2439 = 9'h103 == r_count_5_io_out ? io_r_259_b : _GEN_2438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2440 = 9'h104 == r_count_5_io_out ? io_r_260_b : _GEN_2439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2441 = 9'h105 == r_count_5_io_out ? io_r_261_b : _GEN_2440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2442 = 9'h106 == r_count_5_io_out ? io_r_262_b : _GEN_2441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2443 = 9'h107 == r_count_5_io_out ? io_r_263_b : _GEN_2442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2444 = 9'h108 == r_count_5_io_out ? io_r_264_b : _GEN_2443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2445 = 9'h109 == r_count_5_io_out ? io_r_265_b : _GEN_2444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2446 = 9'h10a == r_count_5_io_out ? io_r_266_b : _GEN_2445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2447 = 9'h10b == r_count_5_io_out ? io_r_267_b : _GEN_2446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2448 = 9'h10c == r_count_5_io_out ? io_r_268_b : _GEN_2447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2449 = 9'h10d == r_count_5_io_out ? io_r_269_b : _GEN_2448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2450 = 9'h10e == r_count_5_io_out ? io_r_270_b : _GEN_2449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2451 = 9'h10f == r_count_5_io_out ? io_r_271_b : _GEN_2450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2452 = 9'h110 == r_count_5_io_out ? io_r_272_b : _GEN_2451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2453 = 9'h111 == r_count_5_io_out ? io_r_273_b : _GEN_2452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2454 = 9'h112 == r_count_5_io_out ? io_r_274_b : _GEN_2453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2455 = 9'h113 == r_count_5_io_out ? io_r_275_b : _GEN_2454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2456 = 9'h114 == r_count_5_io_out ? io_r_276_b : _GEN_2455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2457 = 9'h115 == r_count_5_io_out ? io_r_277_b : _GEN_2456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2458 = 9'h116 == r_count_5_io_out ? io_r_278_b : _GEN_2457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2459 = 9'h117 == r_count_5_io_out ? io_r_279_b : _GEN_2458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2460 = 9'h118 == r_count_5_io_out ? io_r_280_b : _GEN_2459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2461 = 9'h119 == r_count_5_io_out ? io_r_281_b : _GEN_2460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2462 = 9'h11a == r_count_5_io_out ? io_r_282_b : _GEN_2461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2463 = 9'h11b == r_count_5_io_out ? io_r_283_b : _GEN_2462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2464 = 9'h11c == r_count_5_io_out ? io_r_284_b : _GEN_2463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2465 = 9'h11d == r_count_5_io_out ? io_r_285_b : _GEN_2464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2466 = 9'h11e == r_count_5_io_out ? io_r_286_b : _GEN_2465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2467 = 9'h11f == r_count_5_io_out ? io_r_287_b : _GEN_2466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2468 = 9'h120 == r_count_5_io_out ? io_r_288_b : _GEN_2467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2469 = 9'h121 == r_count_5_io_out ? io_r_289_b : _GEN_2468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2470 = 9'h122 == r_count_5_io_out ? io_r_290_b : _GEN_2469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2471 = 9'h123 == r_count_5_io_out ? io_r_291_b : _GEN_2470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2472 = 9'h124 == r_count_5_io_out ? io_r_292_b : _GEN_2471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2473 = 9'h125 == r_count_5_io_out ? io_r_293_b : _GEN_2472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2474 = 9'h126 == r_count_5_io_out ? io_r_294_b : _GEN_2473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2475 = 9'h127 == r_count_5_io_out ? io_r_295_b : _GEN_2474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2476 = 9'h128 == r_count_5_io_out ? io_r_296_b : _GEN_2475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2477 = 9'h129 == r_count_5_io_out ? io_r_297_b : _GEN_2476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2478 = 9'h12a == r_count_5_io_out ? io_r_298_b : _GEN_2477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2479 = 9'h12b == r_count_5_io_out ? io_r_299_b : _GEN_2478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2480 = 9'h12c == r_count_5_io_out ? io_r_300_b : _GEN_2479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2481 = 9'h12d == r_count_5_io_out ? io_r_301_b : _GEN_2480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2482 = 9'h12e == r_count_5_io_out ? io_r_302_b : _GEN_2481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2483 = 9'h12f == r_count_5_io_out ? io_r_303_b : _GEN_2482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2484 = 9'h130 == r_count_5_io_out ? io_r_304_b : _GEN_2483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2485 = 9'h131 == r_count_5_io_out ? io_r_305_b : _GEN_2484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2486 = 9'h132 == r_count_5_io_out ? io_r_306_b : _GEN_2485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2487 = 9'h133 == r_count_5_io_out ? io_r_307_b : _GEN_2486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2488 = 9'h134 == r_count_5_io_out ? io_r_308_b : _GEN_2487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2489 = 9'h135 == r_count_5_io_out ? io_r_309_b : _GEN_2488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2490 = 9'h136 == r_count_5_io_out ? io_r_310_b : _GEN_2489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2491 = 9'h137 == r_count_5_io_out ? io_r_311_b : _GEN_2490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2492 = 9'h138 == r_count_5_io_out ? io_r_312_b : _GEN_2491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2493 = 9'h139 == r_count_5_io_out ? io_r_313_b : _GEN_2492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2494 = 9'h13a == r_count_5_io_out ? io_r_314_b : _GEN_2493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2495 = 9'h13b == r_count_5_io_out ? io_r_315_b : _GEN_2494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2496 = 9'h13c == r_count_5_io_out ? io_r_316_b : _GEN_2495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2497 = 9'h13d == r_count_5_io_out ? io_r_317_b : _GEN_2496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2498 = 9'h13e == r_count_5_io_out ? io_r_318_b : _GEN_2497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2499 = 9'h13f == r_count_5_io_out ? io_r_319_b : _GEN_2498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2500 = 9'h140 == r_count_5_io_out ? io_r_320_b : _GEN_2499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2501 = 9'h141 == r_count_5_io_out ? io_r_321_b : _GEN_2500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2502 = 9'h142 == r_count_5_io_out ? io_r_322_b : _GEN_2501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2503 = 9'h143 == r_count_5_io_out ? io_r_323_b : _GEN_2502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2504 = 9'h144 == r_count_5_io_out ? io_r_324_b : _GEN_2503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2505 = 9'h145 == r_count_5_io_out ? io_r_325_b : _GEN_2504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2506 = 9'h146 == r_count_5_io_out ? io_r_326_b : _GEN_2505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2507 = 9'h147 == r_count_5_io_out ? io_r_327_b : _GEN_2506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2508 = 9'h148 == r_count_5_io_out ? io_r_328_b : _GEN_2507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2509 = 9'h149 == r_count_5_io_out ? io_r_329_b : _GEN_2508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2510 = 9'h14a == r_count_5_io_out ? io_r_330_b : _GEN_2509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2511 = 9'h14b == r_count_5_io_out ? io_r_331_b : _GEN_2510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2512 = 9'h14c == r_count_5_io_out ? io_r_332_b : _GEN_2511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2513 = 9'h14d == r_count_5_io_out ? io_r_333_b : _GEN_2512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2514 = 9'h14e == r_count_5_io_out ? io_r_334_b : _GEN_2513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2515 = 9'h14f == r_count_5_io_out ? io_r_335_b : _GEN_2514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2516 = 9'h150 == r_count_5_io_out ? io_r_336_b : _GEN_2515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2517 = 9'h151 == r_count_5_io_out ? io_r_337_b : _GEN_2516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2518 = 9'h152 == r_count_5_io_out ? io_r_338_b : _GEN_2517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2519 = 9'h153 == r_count_5_io_out ? io_r_339_b : _GEN_2518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2520 = 9'h154 == r_count_5_io_out ? io_r_340_b : _GEN_2519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2521 = 9'h155 == r_count_5_io_out ? io_r_341_b : _GEN_2520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2522 = 9'h156 == r_count_5_io_out ? io_r_342_b : _GEN_2521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2523 = 9'h157 == r_count_5_io_out ? io_r_343_b : _GEN_2522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2524 = 9'h158 == r_count_5_io_out ? io_r_344_b : _GEN_2523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2525 = 9'h159 == r_count_5_io_out ? io_r_345_b : _GEN_2524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2526 = 9'h15a == r_count_5_io_out ? io_r_346_b : _GEN_2525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2527 = 9'h15b == r_count_5_io_out ? io_r_347_b : _GEN_2526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2528 = 9'h15c == r_count_5_io_out ? io_r_348_b : _GEN_2527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2529 = 9'h15d == r_count_5_io_out ? io_r_349_b : _GEN_2528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2530 = 9'h15e == r_count_5_io_out ? io_r_350_b : _GEN_2529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2531 = 9'h15f == r_count_5_io_out ? io_r_351_b : _GEN_2530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2532 = 9'h160 == r_count_5_io_out ? io_r_352_b : _GEN_2531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2533 = 9'h161 == r_count_5_io_out ? io_r_353_b : _GEN_2532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2534 = 9'h162 == r_count_5_io_out ? io_r_354_b : _GEN_2533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2535 = 9'h163 == r_count_5_io_out ? io_r_355_b : _GEN_2534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2536 = 9'h164 == r_count_5_io_out ? io_r_356_b : _GEN_2535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2537 = 9'h165 == r_count_5_io_out ? io_r_357_b : _GEN_2536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2538 = 9'h166 == r_count_5_io_out ? io_r_358_b : _GEN_2537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2539 = 9'h167 == r_count_5_io_out ? io_r_359_b : _GEN_2538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2540 = 9'h168 == r_count_5_io_out ? io_r_360_b : _GEN_2539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2541 = 9'h169 == r_count_5_io_out ? io_r_361_b : _GEN_2540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2542 = 9'h16a == r_count_5_io_out ? io_r_362_b : _GEN_2541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2543 = 9'h16b == r_count_5_io_out ? io_r_363_b : _GEN_2542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2544 = 9'h16c == r_count_5_io_out ? io_r_364_b : _GEN_2543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2545 = 9'h16d == r_count_5_io_out ? io_r_365_b : _GEN_2544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2546 = 9'h16e == r_count_5_io_out ? io_r_366_b : _GEN_2545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2547 = 9'h16f == r_count_5_io_out ? io_r_367_b : _GEN_2546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2548 = 9'h170 == r_count_5_io_out ? io_r_368_b : _GEN_2547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2549 = 9'h171 == r_count_5_io_out ? io_r_369_b : _GEN_2548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2550 = 9'h172 == r_count_5_io_out ? io_r_370_b : _GEN_2549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2551 = 9'h173 == r_count_5_io_out ? io_r_371_b : _GEN_2550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2552 = 9'h174 == r_count_5_io_out ? io_r_372_b : _GEN_2551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2553 = 9'h175 == r_count_5_io_out ? io_r_373_b : _GEN_2552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2554 = 9'h176 == r_count_5_io_out ? io_r_374_b : _GEN_2553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2555 = 9'h177 == r_count_5_io_out ? io_r_375_b : _GEN_2554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2556 = 9'h178 == r_count_5_io_out ? io_r_376_b : _GEN_2555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2557 = 9'h179 == r_count_5_io_out ? io_r_377_b : _GEN_2556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2558 = 9'h17a == r_count_5_io_out ? io_r_378_b : _GEN_2557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2559 = 9'h17b == r_count_5_io_out ? io_r_379_b : _GEN_2558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2560 = 9'h17c == r_count_5_io_out ? io_r_380_b : _GEN_2559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2561 = 9'h17d == r_count_5_io_out ? io_r_381_b : _GEN_2560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2562 = 9'h17e == r_count_5_io_out ? io_r_382_b : _GEN_2561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2563 = 9'h17f == r_count_5_io_out ? io_r_383_b : _GEN_2562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2564 = 9'h180 == r_count_5_io_out ? io_r_384_b : _GEN_2563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2565 = 9'h181 == r_count_5_io_out ? io_r_385_b : _GEN_2564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2566 = 9'h182 == r_count_5_io_out ? io_r_386_b : _GEN_2565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2567 = 9'h183 == r_count_5_io_out ? io_r_387_b : _GEN_2566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2568 = 9'h184 == r_count_5_io_out ? io_r_388_b : _GEN_2567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2569 = 9'h185 == r_count_5_io_out ? io_r_389_b : _GEN_2568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2570 = 9'h186 == r_count_5_io_out ? io_r_390_b : _GEN_2569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2571 = 9'h187 == r_count_5_io_out ? io_r_391_b : _GEN_2570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2572 = 9'h188 == r_count_5_io_out ? io_r_392_b : _GEN_2571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2573 = 9'h189 == r_count_5_io_out ? io_r_393_b : _GEN_2572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2574 = 9'h18a == r_count_5_io_out ? io_r_394_b : _GEN_2573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2575 = 9'h18b == r_count_5_io_out ? io_r_395_b : _GEN_2574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2576 = 9'h18c == r_count_5_io_out ? io_r_396_b : _GEN_2575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2577 = 9'h18d == r_count_5_io_out ? io_r_397_b : _GEN_2576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2578 = 9'h18e == r_count_5_io_out ? io_r_398_b : _GEN_2577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2581 = 9'h1 == r_count_6_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2582 = 9'h2 == r_count_6_io_out ? io_r_2_b : _GEN_2581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2583 = 9'h3 == r_count_6_io_out ? io_r_3_b : _GEN_2582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2584 = 9'h4 == r_count_6_io_out ? io_r_4_b : _GEN_2583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2585 = 9'h5 == r_count_6_io_out ? io_r_5_b : _GEN_2584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2586 = 9'h6 == r_count_6_io_out ? io_r_6_b : _GEN_2585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2587 = 9'h7 == r_count_6_io_out ? io_r_7_b : _GEN_2586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2588 = 9'h8 == r_count_6_io_out ? io_r_8_b : _GEN_2587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2589 = 9'h9 == r_count_6_io_out ? io_r_9_b : _GEN_2588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2590 = 9'ha == r_count_6_io_out ? io_r_10_b : _GEN_2589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2591 = 9'hb == r_count_6_io_out ? io_r_11_b : _GEN_2590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2592 = 9'hc == r_count_6_io_out ? io_r_12_b : _GEN_2591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2593 = 9'hd == r_count_6_io_out ? io_r_13_b : _GEN_2592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2594 = 9'he == r_count_6_io_out ? io_r_14_b : _GEN_2593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2595 = 9'hf == r_count_6_io_out ? io_r_15_b : _GEN_2594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2596 = 9'h10 == r_count_6_io_out ? io_r_16_b : _GEN_2595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2597 = 9'h11 == r_count_6_io_out ? io_r_17_b : _GEN_2596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2598 = 9'h12 == r_count_6_io_out ? io_r_18_b : _GEN_2597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2599 = 9'h13 == r_count_6_io_out ? io_r_19_b : _GEN_2598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2600 = 9'h14 == r_count_6_io_out ? io_r_20_b : _GEN_2599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2601 = 9'h15 == r_count_6_io_out ? io_r_21_b : _GEN_2600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2602 = 9'h16 == r_count_6_io_out ? io_r_22_b : _GEN_2601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2603 = 9'h17 == r_count_6_io_out ? io_r_23_b : _GEN_2602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2604 = 9'h18 == r_count_6_io_out ? io_r_24_b : _GEN_2603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2605 = 9'h19 == r_count_6_io_out ? io_r_25_b : _GEN_2604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2606 = 9'h1a == r_count_6_io_out ? io_r_26_b : _GEN_2605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2607 = 9'h1b == r_count_6_io_out ? io_r_27_b : _GEN_2606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2608 = 9'h1c == r_count_6_io_out ? io_r_28_b : _GEN_2607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2609 = 9'h1d == r_count_6_io_out ? io_r_29_b : _GEN_2608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2610 = 9'h1e == r_count_6_io_out ? io_r_30_b : _GEN_2609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2611 = 9'h1f == r_count_6_io_out ? io_r_31_b : _GEN_2610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2612 = 9'h20 == r_count_6_io_out ? io_r_32_b : _GEN_2611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2613 = 9'h21 == r_count_6_io_out ? io_r_33_b : _GEN_2612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2614 = 9'h22 == r_count_6_io_out ? io_r_34_b : _GEN_2613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2615 = 9'h23 == r_count_6_io_out ? io_r_35_b : _GEN_2614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2616 = 9'h24 == r_count_6_io_out ? io_r_36_b : _GEN_2615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2617 = 9'h25 == r_count_6_io_out ? io_r_37_b : _GEN_2616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2618 = 9'h26 == r_count_6_io_out ? io_r_38_b : _GEN_2617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2619 = 9'h27 == r_count_6_io_out ? io_r_39_b : _GEN_2618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2620 = 9'h28 == r_count_6_io_out ? io_r_40_b : _GEN_2619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2621 = 9'h29 == r_count_6_io_out ? io_r_41_b : _GEN_2620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2622 = 9'h2a == r_count_6_io_out ? io_r_42_b : _GEN_2621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2623 = 9'h2b == r_count_6_io_out ? io_r_43_b : _GEN_2622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2624 = 9'h2c == r_count_6_io_out ? io_r_44_b : _GEN_2623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2625 = 9'h2d == r_count_6_io_out ? io_r_45_b : _GEN_2624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2626 = 9'h2e == r_count_6_io_out ? io_r_46_b : _GEN_2625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2627 = 9'h2f == r_count_6_io_out ? io_r_47_b : _GEN_2626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2628 = 9'h30 == r_count_6_io_out ? io_r_48_b : _GEN_2627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2629 = 9'h31 == r_count_6_io_out ? io_r_49_b : _GEN_2628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2630 = 9'h32 == r_count_6_io_out ? io_r_50_b : _GEN_2629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2631 = 9'h33 == r_count_6_io_out ? io_r_51_b : _GEN_2630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2632 = 9'h34 == r_count_6_io_out ? io_r_52_b : _GEN_2631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2633 = 9'h35 == r_count_6_io_out ? io_r_53_b : _GEN_2632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2634 = 9'h36 == r_count_6_io_out ? io_r_54_b : _GEN_2633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2635 = 9'h37 == r_count_6_io_out ? io_r_55_b : _GEN_2634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2636 = 9'h38 == r_count_6_io_out ? io_r_56_b : _GEN_2635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2637 = 9'h39 == r_count_6_io_out ? io_r_57_b : _GEN_2636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2638 = 9'h3a == r_count_6_io_out ? io_r_58_b : _GEN_2637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2639 = 9'h3b == r_count_6_io_out ? io_r_59_b : _GEN_2638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2640 = 9'h3c == r_count_6_io_out ? io_r_60_b : _GEN_2639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2641 = 9'h3d == r_count_6_io_out ? io_r_61_b : _GEN_2640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2642 = 9'h3e == r_count_6_io_out ? io_r_62_b : _GEN_2641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2643 = 9'h3f == r_count_6_io_out ? io_r_63_b : _GEN_2642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2644 = 9'h40 == r_count_6_io_out ? io_r_64_b : _GEN_2643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2645 = 9'h41 == r_count_6_io_out ? io_r_65_b : _GEN_2644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2646 = 9'h42 == r_count_6_io_out ? io_r_66_b : _GEN_2645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2647 = 9'h43 == r_count_6_io_out ? io_r_67_b : _GEN_2646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2648 = 9'h44 == r_count_6_io_out ? io_r_68_b : _GEN_2647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2649 = 9'h45 == r_count_6_io_out ? io_r_69_b : _GEN_2648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2650 = 9'h46 == r_count_6_io_out ? io_r_70_b : _GEN_2649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2651 = 9'h47 == r_count_6_io_out ? io_r_71_b : _GEN_2650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2652 = 9'h48 == r_count_6_io_out ? io_r_72_b : _GEN_2651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2653 = 9'h49 == r_count_6_io_out ? io_r_73_b : _GEN_2652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2654 = 9'h4a == r_count_6_io_out ? io_r_74_b : _GEN_2653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2655 = 9'h4b == r_count_6_io_out ? io_r_75_b : _GEN_2654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2656 = 9'h4c == r_count_6_io_out ? io_r_76_b : _GEN_2655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2657 = 9'h4d == r_count_6_io_out ? io_r_77_b : _GEN_2656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2658 = 9'h4e == r_count_6_io_out ? io_r_78_b : _GEN_2657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2659 = 9'h4f == r_count_6_io_out ? io_r_79_b : _GEN_2658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2660 = 9'h50 == r_count_6_io_out ? io_r_80_b : _GEN_2659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2661 = 9'h51 == r_count_6_io_out ? io_r_81_b : _GEN_2660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2662 = 9'h52 == r_count_6_io_out ? io_r_82_b : _GEN_2661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2663 = 9'h53 == r_count_6_io_out ? io_r_83_b : _GEN_2662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2664 = 9'h54 == r_count_6_io_out ? io_r_84_b : _GEN_2663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2665 = 9'h55 == r_count_6_io_out ? io_r_85_b : _GEN_2664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2666 = 9'h56 == r_count_6_io_out ? io_r_86_b : _GEN_2665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2667 = 9'h57 == r_count_6_io_out ? io_r_87_b : _GEN_2666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2668 = 9'h58 == r_count_6_io_out ? io_r_88_b : _GEN_2667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2669 = 9'h59 == r_count_6_io_out ? io_r_89_b : _GEN_2668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2670 = 9'h5a == r_count_6_io_out ? io_r_90_b : _GEN_2669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2671 = 9'h5b == r_count_6_io_out ? io_r_91_b : _GEN_2670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2672 = 9'h5c == r_count_6_io_out ? io_r_92_b : _GEN_2671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2673 = 9'h5d == r_count_6_io_out ? io_r_93_b : _GEN_2672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2674 = 9'h5e == r_count_6_io_out ? io_r_94_b : _GEN_2673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2675 = 9'h5f == r_count_6_io_out ? io_r_95_b : _GEN_2674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2676 = 9'h60 == r_count_6_io_out ? io_r_96_b : _GEN_2675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2677 = 9'h61 == r_count_6_io_out ? io_r_97_b : _GEN_2676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2678 = 9'h62 == r_count_6_io_out ? io_r_98_b : _GEN_2677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2679 = 9'h63 == r_count_6_io_out ? io_r_99_b : _GEN_2678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2680 = 9'h64 == r_count_6_io_out ? io_r_100_b : _GEN_2679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2681 = 9'h65 == r_count_6_io_out ? io_r_101_b : _GEN_2680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2682 = 9'h66 == r_count_6_io_out ? io_r_102_b : _GEN_2681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2683 = 9'h67 == r_count_6_io_out ? io_r_103_b : _GEN_2682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2684 = 9'h68 == r_count_6_io_out ? io_r_104_b : _GEN_2683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2685 = 9'h69 == r_count_6_io_out ? io_r_105_b : _GEN_2684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2686 = 9'h6a == r_count_6_io_out ? io_r_106_b : _GEN_2685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2687 = 9'h6b == r_count_6_io_out ? io_r_107_b : _GEN_2686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2688 = 9'h6c == r_count_6_io_out ? io_r_108_b : _GEN_2687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2689 = 9'h6d == r_count_6_io_out ? io_r_109_b : _GEN_2688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2690 = 9'h6e == r_count_6_io_out ? io_r_110_b : _GEN_2689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2691 = 9'h6f == r_count_6_io_out ? io_r_111_b : _GEN_2690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2692 = 9'h70 == r_count_6_io_out ? io_r_112_b : _GEN_2691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2693 = 9'h71 == r_count_6_io_out ? io_r_113_b : _GEN_2692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2694 = 9'h72 == r_count_6_io_out ? io_r_114_b : _GEN_2693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2695 = 9'h73 == r_count_6_io_out ? io_r_115_b : _GEN_2694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2696 = 9'h74 == r_count_6_io_out ? io_r_116_b : _GEN_2695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2697 = 9'h75 == r_count_6_io_out ? io_r_117_b : _GEN_2696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2698 = 9'h76 == r_count_6_io_out ? io_r_118_b : _GEN_2697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2699 = 9'h77 == r_count_6_io_out ? io_r_119_b : _GEN_2698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2700 = 9'h78 == r_count_6_io_out ? io_r_120_b : _GEN_2699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2701 = 9'h79 == r_count_6_io_out ? io_r_121_b : _GEN_2700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2702 = 9'h7a == r_count_6_io_out ? io_r_122_b : _GEN_2701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2703 = 9'h7b == r_count_6_io_out ? io_r_123_b : _GEN_2702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2704 = 9'h7c == r_count_6_io_out ? io_r_124_b : _GEN_2703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2705 = 9'h7d == r_count_6_io_out ? io_r_125_b : _GEN_2704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2706 = 9'h7e == r_count_6_io_out ? io_r_126_b : _GEN_2705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2707 = 9'h7f == r_count_6_io_out ? io_r_127_b : _GEN_2706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2708 = 9'h80 == r_count_6_io_out ? io_r_128_b : _GEN_2707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2709 = 9'h81 == r_count_6_io_out ? io_r_129_b : _GEN_2708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2710 = 9'h82 == r_count_6_io_out ? io_r_130_b : _GEN_2709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2711 = 9'h83 == r_count_6_io_out ? io_r_131_b : _GEN_2710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2712 = 9'h84 == r_count_6_io_out ? io_r_132_b : _GEN_2711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2713 = 9'h85 == r_count_6_io_out ? io_r_133_b : _GEN_2712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2714 = 9'h86 == r_count_6_io_out ? io_r_134_b : _GEN_2713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2715 = 9'h87 == r_count_6_io_out ? io_r_135_b : _GEN_2714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2716 = 9'h88 == r_count_6_io_out ? io_r_136_b : _GEN_2715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2717 = 9'h89 == r_count_6_io_out ? io_r_137_b : _GEN_2716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2718 = 9'h8a == r_count_6_io_out ? io_r_138_b : _GEN_2717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2719 = 9'h8b == r_count_6_io_out ? io_r_139_b : _GEN_2718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2720 = 9'h8c == r_count_6_io_out ? io_r_140_b : _GEN_2719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2721 = 9'h8d == r_count_6_io_out ? io_r_141_b : _GEN_2720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2722 = 9'h8e == r_count_6_io_out ? io_r_142_b : _GEN_2721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2723 = 9'h8f == r_count_6_io_out ? io_r_143_b : _GEN_2722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2724 = 9'h90 == r_count_6_io_out ? io_r_144_b : _GEN_2723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2725 = 9'h91 == r_count_6_io_out ? io_r_145_b : _GEN_2724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2726 = 9'h92 == r_count_6_io_out ? io_r_146_b : _GEN_2725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2727 = 9'h93 == r_count_6_io_out ? io_r_147_b : _GEN_2726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2728 = 9'h94 == r_count_6_io_out ? io_r_148_b : _GEN_2727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2729 = 9'h95 == r_count_6_io_out ? io_r_149_b : _GEN_2728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2730 = 9'h96 == r_count_6_io_out ? io_r_150_b : _GEN_2729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2731 = 9'h97 == r_count_6_io_out ? io_r_151_b : _GEN_2730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2732 = 9'h98 == r_count_6_io_out ? io_r_152_b : _GEN_2731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2733 = 9'h99 == r_count_6_io_out ? io_r_153_b : _GEN_2732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2734 = 9'h9a == r_count_6_io_out ? io_r_154_b : _GEN_2733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2735 = 9'h9b == r_count_6_io_out ? io_r_155_b : _GEN_2734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2736 = 9'h9c == r_count_6_io_out ? io_r_156_b : _GEN_2735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2737 = 9'h9d == r_count_6_io_out ? io_r_157_b : _GEN_2736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2738 = 9'h9e == r_count_6_io_out ? io_r_158_b : _GEN_2737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2739 = 9'h9f == r_count_6_io_out ? io_r_159_b : _GEN_2738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2740 = 9'ha0 == r_count_6_io_out ? io_r_160_b : _GEN_2739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2741 = 9'ha1 == r_count_6_io_out ? io_r_161_b : _GEN_2740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2742 = 9'ha2 == r_count_6_io_out ? io_r_162_b : _GEN_2741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2743 = 9'ha3 == r_count_6_io_out ? io_r_163_b : _GEN_2742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2744 = 9'ha4 == r_count_6_io_out ? io_r_164_b : _GEN_2743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2745 = 9'ha5 == r_count_6_io_out ? io_r_165_b : _GEN_2744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2746 = 9'ha6 == r_count_6_io_out ? io_r_166_b : _GEN_2745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2747 = 9'ha7 == r_count_6_io_out ? io_r_167_b : _GEN_2746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2748 = 9'ha8 == r_count_6_io_out ? io_r_168_b : _GEN_2747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2749 = 9'ha9 == r_count_6_io_out ? io_r_169_b : _GEN_2748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2750 = 9'haa == r_count_6_io_out ? io_r_170_b : _GEN_2749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2751 = 9'hab == r_count_6_io_out ? io_r_171_b : _GEN_2750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2752 = 9'hac == r_count_6_io_out ? io_r_172_b : _GEN_2751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2753 = 9'had == r_count_6_io_out ? io_r_173_b : _GEN_2752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2754 = 9'hae == r_count_6_io_out ? io_r_174_b : _GEN_2753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2755 = 9'haf == r_count_6_io_out ? io_r_175_b : _GEN_2754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2756 = 9'hb0 == r_count_6_io_out ? io_r_176_b : _GEN_2755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2757 = 9'hb1 == r_count_6_io_out ? io_r_177_b : _GEN_2756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2758 = 9'hb2 == r_count_6_io_out ? io_r_178_b : _GEN_2757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2759 = 9'hb3 == r_count_6_io_out ? io_r_179_b : _GEN_2758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2760 = 9'hb4 == r_count_6_io_out ? io_r_180_b : _GEN_2759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2761 = 9'hb5 == r_count_6_io_out ? io_r_181_b : _GEN_2760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2762 = 9'hb6 == r_count_6_io_out ? io_r_182_b : _GEN_2761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2763 = 9'hb7 == r_count_6_io_out ? io_r_183_b : _GEN_2762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2764 = 9'hb8 == r_count_6_io_out ? io_r_184_b : _GEN_2763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2765 = 9'hb9 == r_count_6_io_out ? io_r_185_b : _GEN_2764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2766 = 9'hba == r_count_6_io_out ? io_r_186_b : _GEN_2765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2767 = 9'hbb == r_count_6_io_out ? io_r_187_b : _GEN_2766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2768 = 9'hbc == r_count_6_io_out ? io_r_188_b : _GEN_2767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2769 = 9'hbd == r_count_6_io_out ? io_r_189_b : _GEN_2768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2770 = 9'hbe == r_count_6_io_out ? io_r_190_b : _GEN_2769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2771 = 9'hbf == r_count_6_io_out ? io_r_191_b : _GEN_2770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2772 = 9'hc0 == r_count_6_io_out ? io_r_192_b : _GEN_2771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2773 = 9'hc1 == r_count_6_io_out ? io_r_193_b : _GEN_2772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2774 = 9'hc2 == r_count_6_io_out ? io_r_194_b : _GEN_2773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2775 = 9'hc3 == r_count_6_io_out ? io_r_195_b : _GEN_2774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2776 = 9'hc4 == r_count_6_io_out ? io_r_196_b : _GEN_2775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2777 = 9'hc5 == r_count_6_io_out ? io_r_197_b : _GEN_2776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2778 = 9'hc6 == r_count_6_io_out ? io_r_198_b : _GEN_2777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2779 = 9'hc7 == r_count_6_io_out ? io_r_199_b : _GEN_2778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2780 = 9'hc8 == r_count_6_io_out ? io_r_200_b : _GEN_2779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2781 = 9'hc9 == r_count_6_io_out ? io_r_201_b : _GEN_2780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2782 = 9'hca == r_count_6_io_out ? io_r_202_b : _GEN_2781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2783 = 9'hcb == r_count_6_io_out ? io_r_203_b : _GEN_2782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2784 = 9'hcc == r_count_6_io_out ? io_r_204_b : _GEN_2783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2785 = 9'hcd == r_count_6_io_out ? io_r_205_b : _GEN_2784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2786 = 9'hce == r_count_6_io_out ? io_r_206_b : _GEN_2785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2787 = 9'hcf == r_count_6_io_out ? io_r_207_b : _GEN_2786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2788 = 9'hd0 == r_count_6_io_out ? io_r_208_b : _GEN_2787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2789 = 9'hd1 == r_count_6_io_out ? io_r_209_b : _GEN_2788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2790 = 9'hd2 == r_count_6_io_out ? io_r_210_b : _GEN_2789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2791 = 9'hd3 == r_count_6_io_out ? io_r_211_b : _GEN_2790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2792 = 9'hd4 == r_count_6_io_out ? io_r_212_b : _GEN_2791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2793 = 9'hd5 == r_count_6_io_out ? io_r_213_b : _GEN_2792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2794 = 9'hd6 == r_count_6_io_out ? io_r_214_b : _GEN_2793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2795 = 9'hd7 == r_count_6_io_out ? io_r_215_b : _GEN_2794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2796 = 9'hd8 == r_count_6_io_out ? io_r_216_b : _GEN_2795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2797 = 9'hd9 == r_count_6_io_out ? io_r_217_b : _GEN_2796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2798 = 9'hda == r_count_6_io_out ? io_r_218_b : _GEN_2797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2799 = 9'hdb == r_count_6_io_out ? io_r_219_b : _GEN_2798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2800 = 9'hdc == r_count_6_io_out ? io_r_220_b : _GEN_2799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2801 = 9'hdd == r_count_6_io_out ? io_r_221_b : _GEN_2800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2802 = 9'hde == r_count_6_io_out ? io_r_222_b : _GEN_2801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2803 = 9'hdf == r_count_6_io_out ? io_r_223_b : _GEN_2802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2804 = 9'he0 == r_count_6_io_out ? io_r_224_b : _GEN_2803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2805 = 9'he1 == r_count_6_io_out ? io_r_225_b : _GEN_2804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2806 = 9'he2 == r_count_6_io_out ? io_r_226_b : _GEN_2805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2807 = 9'he3 == r_count_6_io_out ? io_r_227_b : _GEN_2806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2808 = 9'he4 == r_count_6_io_out ? io_r_228_b : _GEN_2807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2809 = 9'he5 == r_count_6_io_out ? io_r_229_b : _GEN_2808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2810 = 9'he6 == r_count_6_io_out ? io_r_230_b : _GEN_2809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2811 = 9'he7 == r_count_6_io_out ? io_r_231_b : _GEN_2810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2812 = 9'he8 == r_count_6_io_out ? io_r_232_b : _GEN_2811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2813 = 9'he9 == r_count_6_io_out ? io_r_233_b : _GEN_2812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2814 = 9'hea == r_count_6_io_out ? io_r_234_b : _GEN_2813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2815 = 9'heb == r_count_6_io_out ? io_r_235_b : _GEN_2814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2816 = 9'hec == r_count_6_io_out ? io_r_236_b : _GEN_2815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2817 = 9'hed == r_count_6_io_out ? io_r_237_b : _GEN_2816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2818 = 9'hee == r_count_6_io_out ? io_r_238_b : _GEN_2817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2819 = 9'hef == r_count_6_io_out ? io_r_239_b : _GEN_2818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2820 = 9'hf0 == r_count_6_io_out ? io_r_240_b : _GEN_2819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2821 = 9'hf1 == r_count_6_io_out ? io_r_241_b : _GEN_2820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2822 = 9'hf2 == r_count_6_io_out ? io_r_242_b : _GEN_2821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2823 = 9'hf3 == r_count_6_io_out ? io_r_243_b : _GEN_2822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2824 = 9'hf4 == r_count_6_io_out ? io_r_244_b : _GEN_2823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2825 = 9'hf5 == r_count_6_io_out ? io_r_245_b : _GEN_2824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2826 = 9'hf6 == r_count_6_io_out ? io_r_246_b : _GEN_2825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2827 = 9'hf7 == r_count_6_io_out ? io_r_247_b : _GEN_2826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2828 = 9'hf8 == r_count_6_io_out ? io_r_248_b : _GEN_2827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2829 = 9'hf9 == r_count_6_io_out ? io_r_249_b : _GEN_2828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2830 = 9'hfa == r_count_6_io_out ? io_r_250_b : _GEN_2829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2831 = 9'hfb == r_count_6_io_out ? io_r_251_b : _GEN_2830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2832 = 9'hfc == r_count_6_io_out ? io_r_252_b : _GEN_2831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2833 = 9'hfd == r_count_6_io_out ? io_r_253_b : _GEN_2832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2834 = 9'hfe == r_count_6_io_out ? io_r_254_b : _GEN_2833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2835 = 9'hff == r_count_6_io_out ? io_r_255_b : _GEN_2834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2836 = 9'h100 == r_count_6_io_out ? io_r_256_b : _GEN_2835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2837 = 9'h101 == r_count_6_io_out ? io_r_257_b : _GEN_2836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2838 = 9'h102 == r_count_6_io_out ? io_r_258_b : _GEN_2837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2839 = 9'h103 == r_count_6_io_out ? io_r_259_b : _GEN_2838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2840 = 9'h104 == r_count_6_io_out ? io_r_260_b : _GEN_2839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2841 = 9'h105 == r_count_6_io_out ? io_r_261_b : _GEN_2840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2842 = 9'h106 == r_count_6_io_out ? io_r_262_b : _GEN_2841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2843 = 9'h107 == r_count_6_io_out ? io_r_263_b : _GEN_2842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2844 = 9'h108 == r_count_6_io_out ? io_r_264_b : _GEN_2843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2845 = 9'h109 == r_count_6_io_out ? io_r_265_b : _GEN_2844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2846 = 9'h10a == r_count_6_io_out ? io_r_266_b : _GEN_2845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2847 = 9'h10b == r_count_6_io_out ? io_r_267_b : _GEN_2846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2848 = 9'h10c == r_count_6_io_out ? io_r_268_b : _GEN_2847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2849 = 9'h10d == r_count_6_io_out ? io_r_269_b : _GEN_2848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2850 = 9'h10e == r_count_6_io_out ? io_r_270_b : _GEN_2849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2851 = 9'h10f == r_count_6_io_out ? io_r_271_b : _GEN_2850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2852 = 9'h110 == r_count_6_io_out ? io_r_272_b : _GEN_2851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2853 = 9'h111 == r_count_6_io_out ? io_r_273_b : _GEN_2852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2854 = 9'h112 == r_count_6_io_out ? io_r_274_b : _GEN_2853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2855 = 9'h113 == r_count_6_io_out ? io_r_275_b : _GEN_2854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2856 = 9'h114 == r_count_6_io_out ? io_r_276_b : _GEN_2855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2857 = 9'h115 == r_count_6_io_out ? io_r_277_b : _GEN_2856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2858 = 9'h116 == r_count_6_io_out ? io_r_278_b : _GEN_2857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2859 = 9'h117 == r_count_6_io_out ? io_r_279_b : _GEN_2858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2860 = 9'h118 == r_count_6_io_out ? io_r_280_b : _GEN_2859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2861 = 9'h119 == r_count_6_io_out ? io_r_281_b : _GEN_2860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2862 = 9'h11a == r_count_6_io_out ? io_r_282_b : _GEN_2861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2863 = 9'h11b == r_count_6_io_out ? io_r_283_b : _GEN_2862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2864 = 9'h11c == r_count_6_io_out ? io_r_284_b : _GEN_2863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2865 = 9'h11d == r_count_6_io_out ? io_r_285_b : _GEN_2864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2866 = 9'h11e == r_count_6_io_out ? io_r_286_b : _GEN_2865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2867 = 9'h11f == r_count_6_io_out ? io_r_287_b : _GEN_2866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2868 = 9'h120 == r_count_6_io_out ? io_r_288_b : _GEN_2867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2869 = 9'h121 == r_count_6_io_out ? io_r_289_b : _GEN_2868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2870 = 9'h122 == r_count_6_io_out ? io_r_290_b : _GEN_2869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2871 = 9'h123 == r_count_6_io_out ? io_r_291_b : _GEN_2870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2872 = 9'h124 == r_count_6_io_out ? io_r_292_b : _GEN_2871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2873 = 9'h125 == r_count_6_io_out ? io_r_293_b : _GEN_2872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2874 = 9'h126 == r_count_6_io_out ? io_r_294_b : _GEN_2873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2875 = 9'h127 == r_count_6_io_out ? io_r_295_b : _GEN_2874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2876 = 9'h128 == r_count_6_io_out ? io_r_296_b : _GEN_2875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2877 = 9'h129 == r_count_6_io_out ? io_r_297_b : _GEN_2876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2878 = 9'h12a == r_count_6_io_out ? io_r_298_b : _GEN_2877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2879 = 9'h12b == r_count_6_io_out ? io_r_299_b : _GEN_2878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2880 = 9'h12c == r_count_6_io_out ? io_r_300_b : _GEN_2879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2881 = 9'h12d == r_count_6_io_out ? io_r_301_b : _GEN_2880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2882 = 9'h12e == r_count_6_io_out ? io_r_302_b : _GEN_2881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2883 = 9'h12f == r_count_6_io_out ? io_r_303_b : _GEN_2882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2884 = 9'h130 == r_count_6_io_out ? io_r_304_b : _GEN_2883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2885 = 9'h131 == r_count_6_io_out ? io_r_305_b : _GEN_2884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2886 = 9'h132 == r_count_6_io_out ? io_r_306_b : _GEN_2885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2887 = 9'h133 == r_count_6_io_out ? io_r_307_b : _GEN_2886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2888 = 9'h134 == r_count_6_io_out ? io_r_308_b : _GEN_2887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2889 = 9'h135 == r_count_6_io_out ? io_r_309_b : _GEN_2888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2890 = 9'h136 == r_count_6_io_out ? io_r_310_b : _GEN_2889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2891 = 9'h137 == r_count_6_io_out ? io_r_311_b : _GEN_2890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2892 = 9'h138 == r_count_6_io_out ? io_r_312_b : _GEN_2891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2893 = 9'h139 == r_count_6_io_out ? io_r_313_b : _GEN_2892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2894 = 9'h13a == r_count_6_io_out ? io_r_314_b : _GEN_2893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2895 = 9'h13b == r_count_6_io_out ? io_r_315_b : _GEN_2894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2896 = 9'h13c == r_count_6_io_out ? io_r_316_b : _GEN_2895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2897 = 9'h13d == r_count_6_io_out ? io_r_317_b : _GEN_2896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2898 = 9'h13e == r_count_6_io_out ? io_r_318_b : _GEN_2897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2899 = 9'h13f == r_count_6_io_out ? io_r_319_b : _GEN_2898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2900 = 9'h140 == r_count_6_io_out ? io_r_320_b : _GEN_2899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2901 = 9'h141 == r_count_6_io_out ? io_r_321_b : _GEN_2900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2902 = 9'h142 == r_count_6_io_out ? io_r_322_b : _GEN_2901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2903 = 9'h143 == r_count_6_io_out ? io_r_323_b : _GEN_2902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2904 = 9'h144 == r_count_6_io_out ? io_r_324_b : _GEN_2903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2905 = 9'h145 == r_count_6_io_out ? io_r_325_b : _GEN_2904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2906 = 9'h146 == r_count_6_io_out ? io_r_326_b : _GEN_2905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2907 = 9'h147 == r_count_6_io_out ? io_r_327_b : _GEN_2906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2908 = 9'h148 == r_count_6_io_out ? io_r_328_b : _GEN_2907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2909 = 9'h149 == r_count_6_io_out ? io_r_329_b : _GEN_2908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2910 = 9'h14a == r_count_6_io_out ? io_r_330_b : _GEN_2909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2911 = 9'h14b == r_count_6_io_out ? io_r_331_b : _GEN_2910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2912 = 9'h14c == r_count_6_io_out ? io_r_332_b : _GEN_2911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2913 = 9'h14d == r_count_6_io_out ? io_r_333_b : _GEN_2912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2914 = 9'h14e == r_count_6_io_out ? io_r_334_b : _GEN_2913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2915 = 9'h14f == r_count_6_io_out ? io_r_335_b : _GEN_2914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2916 = 9'h150 == r_count_6_io_out ? io_r_336_b : _GEN_2915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2917 = 9'h151 == r_count_6_io_out ? io_r_337_b : _GEN_2916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2918 = 9'h152 == r_count_6_io_out ? io_r_338_b : _GEN_2917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2919 = 9'h153 == r_count_6_io_out ? io_r_339_b : _GEN_2918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2920 = 9'h154 == r_count_6_io_out ? io_r_340_b : _GEN_2919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2921 = 9'h155 == r_count_6_io_out ? io_r_341_b : _GEN_2920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2922 = 9'h156 == r_count_6_io_out ? io_r_342_b : _GEN_2921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2923 = 9'h157 == r_count_6_io_out ? io_r_343_b : _GEN_2922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2924 = 9'h158 == r_count_6_io_out ? io_r_344_b : _GEN_2923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2925 = 9'h159 == r_count_6_io_out ? io_r_345_b : _GEN_2924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2926 = 9'h15a == r_count_6_io_out ? io_r_346_b : _GEN_2925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2927 = 9'h15b == r_count_6_io_out ? io_r_347_b : _GEN_2926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2928 = 9'h15c == r_count_6_io_out ? io_r_348_b : _GEN_2927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2929 = 9'h15d == r_count_6_io_out ? io_r_349_b : _GEN_2928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2930 = 9'h15e == r_count_6_io_out ? io_r_350_b : _GEN_2929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2931 = 9'h15f == r_count_6_io_out ? io_r_351_b : _GEN_2930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2932 = 9'h160 == r_count_6_io_out ? io_r_352_b : _GEN_2931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2933 = 9'h161 == r_count_6_io_out ? io_r_353_b : _GEN_2932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2934 = 9'h162 == r_count_6_io_out ? io_r_354_b : _GEN_2933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2935 = 9'h163 == r_count_6_io_out ? io_r_355_b : _GEN_2934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2936 = 9'h164 == r_count_6_io_out ? io_r_356_b : _GEN_2935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2937 = 9'h165 == r_count_6_io_out ? io_r_357_b : _GEN_2936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2938 = 9'h166 == r_count_6_io_out ? io_r_358_b : _GEN_2937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2939 = 9'h167 == r_count_6_io_out ? io_r_359_b : _GEN_2938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2940 = 9'h168 == r_count_6_io_out ? io_r_360_b : _GEN_2939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2941 = 9'h169 == r_count_6_io_out ? io_r_361_b : _GEN_2940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2942 = 9'h16a == r_count_6_io_out ? io_r_362_b : _GEN_2941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2943 = 9'h16b == r_count_6_io_out ? io_r_363_b : _GEN_2942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2944 = 9'h16c == r_count_6_io_out ? io_r_364_b : _GEN_2943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2945 = 9'h16d == r_count_6_io_out ? io_r_365_b : _GEN_2944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2946 = 9'h16e == r_count_6_io_out ? io_r_366_b : _GEN_2945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2947 = 9'h16f == r_count_6_io_out ? io_r_367_b : _GEN_2946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2948 = 9'h170 == r_count_6_io_out ? io_r_368_b : _GEN_2947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2949 = 9'h171 == r_count_6_io_out ? io_r_369_b : _GEN_2948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2950 = 9'h172 == r_count_6_io_out ? io_r_370_b : _GEN_2949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2951 = 9'h173 == r_count_6_io_out ? io_r_371_b : _GEN_2950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2952 = 9'h174 == r_count_6_io_out ? io_r_372_b : _GEN_2951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2953 = 9'h175 == r_count_6_io_out ? io_r_373_b : _GEN_2952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2954 = 9'h176 == r_count_6_io_out ? io_r_374_b : _GEN_2953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2955 = 9'h177 == r_count_6_io_out ? io_r_375_b : _GEN_2954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2956 = 9'h178 == r_count_6_io_out ? io_r_376_b : _GEN_2955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2957 = 9'h179 == r_count_6_io_out ? io_r_377_b : _GEN_2956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2958 = 9'h17a == r_count_6_io_out ? io_r_378_b : _GEN_2957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2959 = 9'h17b == r_count_6_io_out ? io_r_379_b : _GEN_2958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2960 = 9'h17c == r_count_6_io_out ? io_r_380_b : _GEN_2959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2961 = 9'h17d == r_count_6_io_out ? io_r_381_b : _GEN_2960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2962 = 9'h17e == r_count_6_io_out ? io_r_382_b : _GEN_2961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2963 = 9'h17f == r_count_6_io_out ? io_r_383_b : _GEN_2962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2964 = 9'h180 == r_count_6_io_out ? io_r_384_b : _GEN_2963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2965 = 9'h181 == r_count_6_io_out ? io_r_385_b : _GEN_2964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2966 = 9'h182 == r_count_6_io_out ? io_r_386_b : _GEN_2965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2967 = 9'h183 == r_count_6_io_out ? io_r_387_b : _GEN_2966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2968 = 9'h184 == r_count_6_io_out ? io_r_388_b : _GEN_2967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2969 = 9'h185 == r_count_6_io_out ? io_r_389_b : _GEN_2968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2970 = 9'h186 == r_count_6_io_out ? io_r_390_b : _GEN_2969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2971 = 9'h187 == r_count_6_io_out ? io_r_391_b : _GEN_2970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2972 = 9'h188 == r_count_6_io_out ? io_r_392_b : _GEN_2971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2973 = 9'h189 == r_count_6_io_out ? io_r_393_b : _GEN_2972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2974 = 9'h18a == r_count_6_io_out ? io_r_394_b : _GEN_2973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2975 = 9'h18b == r_count_6_io_out ? io_r_395_b : _GEN_2974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2976 = 9'h18c == r_count_6_io_out ? io_r_396_b : _GEN_2975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2977 = 9'h18d == r_count_6_io_out ? io_r_397_b : _GEN_2976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2978 = 9'h18e == r_count_6_io_out ? io_r_398_b : _GEN_2977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2981 = 9'h1 == r_count_7_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2982 = 9'h2 == r_count_7_io_out ? io_r_2_b : _GEN_2981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2983 = 9'h3 == r_count_7_io_out ? io_r_3_b : _GEN_2982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2984 = 9'h4 == r_count_7_io_out ? io_r_4_b : _GEN_2983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2985 = 9'h5 == r_count_7_io_out ? io_r_5_b : _GEN_2984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2986 = 9'h6 == r_count_7_io_out ? io_r_6_b : _GEN_2985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2987 = 9'h7 == r_count_7_io_out ? io_r_7_b : _GEN_2986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2988 = 9'h8 == r_count_7_io_out ? io_r_8_b : _GEN_2987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2989 = 9'h9 == r_count_7_io_out ? io_r_9_b : _GEN_2988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2990 = 9'ha == r_count_7_io_out ? io_r_10_b : _GEN_2989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2991 = 9'hb == r_count_7_io_out ? io_r_11_b : _GEN_2990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2992 = 9'hc == r_count_7_io_out ? io_r_12_b : _GEN_2991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2993 = 9'hd == r_count_7_io_out ? io_r_13_b : _GEN_2992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2994 = 9'he == r_count_7_io_out ? io_r_14_b : _GEN_2993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2995 = 9'hf == r_count_7_io_out ? io_r_15_b : _GEN_2994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2996 = 9'h10 == r_count_7_io_out ? io_r_16_b : _GEN_2995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2997 = 9'h11 == r_count_7_io_out ? io_r_17_b : _GEN_2996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2998 = 9'h12 == r_count_7_io_out ? io_r_18_b : _GEN_2997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2999 = 9'h13 == r_count_7_io_out ? io_r_19_b : _GEN_2998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3000 = 9'h14 == r_count_7_io_out ? io_r_20_b : _GEN_2999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3001 = 9'h15 == r_count_7_io_out ? io_r_21_b : _GEN_3000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3002 = 9'h16 == r_count_7_io_out ? io_r_22_b : _GEN_3001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3003 = 9'h17 == r_count_7_io_out ? io_r_23_b : _GEN_3002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3004 = 9'h18 == r_count_7_io_out ? io_r_24_b : _GEN_3003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3005 = 9'h19 == r_count_7_io_out ? io_r_25_b : _GEN_3004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3006 = 9'h1a == r_count_7_io_out ? io_r_26_b : _GEN_3005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3007 = 9'h1b == r_count_7_io_out ? io_r_27_b : _GEN_3006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3008 = 9'h1c == r_count_7_io_out ? io_r_28_b : _GEN_3007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3009 = 9'h1d == r_count_7_io_out ? io_r_29_b : _GEN_3008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3010 = 9'h1e == r_count_7_io_out ? io_r_30_b : _GEN_3009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3011 = 9'h1f == r_count_7_io_out ? io_r_31_b : _GEN_3010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3012 = 9'h20 == r_count_7_io_out ? io_r_32_b : _GEN_3011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3013 = 9'h21 == r_count_7_io_out ? io_r_33_b : _GEN_3012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3014 = 9'h22 == r_count_7_io_out ? io_r_34_b : _GEN_3013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3015 = 9'h23 == r_count_7_io_out ? io_r_35_b : _GEN_3014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3016 = 9'h24 == r_count_7_io_out ? io_r_36_b : _GEN_3015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3017 = 9'h25 == r_count_7_io_out ? io_r_37_b : _GEN_3016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3018 = 9'h26 == r_count_7_io_out ? io_r_38_b : _GEN_3017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3019 = 9'h27 == r_count_7_io_out ? io_r_39_b : _GEN_3018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3020 = 9'h28 == r_count_7_io_out ? io_r_40_b : _GEN_3019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3021 = 9'h29 == r_count_7_io_out ? io_r_41_b : _GEN_3020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3022 = 9'h2a == r_count_7_io_out ? io_r_42_b : _GEN_3021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3023 = 9'h2b == r_count_7_io_out ? io_r_43_b : _GEN_3022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3024 = 9'h2c == r_count_7_io_out ? io_r_44_b : _GEN_3023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3025 = 9'h2d == r_count_7_io_out ? io_r_45_b : _GEN_3024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3026 = 9'h2e == r_count_7_io_out ? io_r_46_b : _GEN_3025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3027 = 9'h2f == r_count_7_io_out ? io_r_47_b : _GEN_3026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3028 = 9'h30 == r_count_7_io_out ? io_r_48_b : _GEN_3027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3029 = 9'h31 == r_count_7_io_out ? io_r_49_b : _GEN_3028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3030 = 9'h32 == r_count_7_io_out ? io_r_50_b : _GEN_3029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3031 = 9'h33 == r_count_7_io_out ? io_r_51_b : _GEN_3030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3032 = 9'h34 == r_count_7_io_out ? io_r_52_b : _GEN_3031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3033 = 9'h35 == r_count_7_io_out ? io_r_53_b : _GEN_3032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3034 = 9'h36 == r_count_7_io_out ? io_r_54_b : _GEN_3033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3035 = 9'h37 == r_count_7_io_out ? io_r_55_b : _GEN_3034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3036 = 9'h38 == r_count_7_io_out ? io_r_56_b : _GEN_3035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3037 = 9'h39 == r_count_7_io_out ? io_r_57_b : _GEN_3036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3038 = 9'h3a == r_count_7_io_out ? io_r_58_b : _GEN_3037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3039 = 9'h3b == r_count_7_io_out ? io_r_59_b : _GEN_3038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3040 = 9'h3c == r_count_7_io_out ? io_r_60_b : _GEN_3039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3041 = 9'h3d == r_count_7_io_out ? io_r_61_b : _GEN_3040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3042 = 9'h3e == r_count_7_io_out ? io_r_62_b : _GEN_3041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3043 = 9'h3f == r_count_7_io_out ? io_r_63_b : _GEN_3042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3044 = 9'h40 == r_count_7_io_out ? io_r_64_b : _GEN_3043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3045 = 9'h41 == r_count_7_io_out ? io_r_65_b : _GEN_3044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3046 = 9'h42 == r_count_7_io_out ? io_r_66_b : _GEN_3045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3047 = 9'h43 == r_count_7_io_out ? io_r_67_b : _GEN_3046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3048 = 9'h44 == r_count_7_io_out ? io_r_68_b : _GEN_3047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3049 = 9'h45 == r_count_7_io_out ? io_r_69_b : _GEN_3048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3050 = 9'h46 == r_count_7_io_out ? io_r_70_b : _GEN_3049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3051 = 9'h47 == r_count_7_io_out ? io_r_71_b : _GEN_3050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3052 = 9'h48 == r_count_7_io_out ? io_r_72_b : _GEN_3051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3053 = 9'h49 == r_count_7_io_out ? io_r_73_b : _GEN_3052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3054 = 9'h4a == r_count_7_io_out ? io_r_74_b : _GEN_3053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3055 = 9'h4b == r_count_7_io_out ? io_r_75_b : _GEN_3054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3056 = 9'h4c == r_count_7_io_out ? io_r_76_b : _GEN_3055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3057 = 9'h4d == r_count_7_io_out ? io_r_77_b : _GEN_3056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3058 = 9'h4e == r_count_7_io_out ? io_r_78_b : _GEN_3057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3059 = 9'h4f == r_count_7_io_out ? io_r_79_b : _GEN_3058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3060 = 9'h50 == r_count_7_io_out ? io_r_80_b : _GEN_3059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3061 = 9'h51 == r_count_7_io_out ? io_r_81_b : _GEN_3060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3062 = 9'h52 == r_count_7_io_out ? io_r_82_b : _GEN_3061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3063 = 9'h53 == r_count_7_io_out ? io_r_83_b : _GEN_3062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3064 = 9'h54 == r_count_7_io_out ? io_r_84_b : _GEN_3063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3065 = 9'h55 == r_count_7_io_out ? io_r_85_b : _GEN_3064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3066 = 9'h56 == r_count_7_io_out ? io_r_86_b : _GEN_3065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3067 = 9'h57 == r_count_7_io_out ? io_r_87_b : _GEN_3066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3068 = 9'h58 == r_count_7_io_out ? io_r_88_b : _GEN_3067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3069 = 9'h59 == r_count_7_io_out ? io_r_89_b : _GEN_3068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3070 = 9'h5a == r_count_7_io_out ? io_r_90_b : _GEN_3069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3071 = 9'h5b == r_count_7_io_out ? io_r_91_b : _GEN_3070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3072 = 9'h5c == r_count_7_io_out ? io_r_92_b : _GEN_3071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3073 = 9'h5d == r_count_7_io_out ? io_r_93_b : _GEN_3072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3074 = 9'h5e == r_count_7_io_out ? io_r_94_b : _GEN_3073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3075 = 9'h5f == r_count_7_io_out ? io_r_95_b : _GEN_3074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3076 = 9'h60 == r_count_7_io_out ? io_r_96_b : _GEN_3075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3077 = 9'h61 == r_count_7_io_out ? io_r_97_b : _GEN_3076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3078 = 9'h62 == r_count_7_io_out ? io_r_98_b : _GEN_3077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3079 = 9'h63 == r_count_7_io_out ? io_r_99_b : _GEN_3078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3080 = 9'h64 == r_count_7_io_out ? io_r_100_b : _GEN_3079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3081 = 9'h65 == r_count_7_io_out ? io_r_101_b : _GEN_3080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3082 = 9'h66 == r_count_7_io_out ? io_r_102_b : _GEN_3081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3083 = 9'h67 == r_count_7_io_out ? io_r_103_b : _GEN_3082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3084 = 9'h68 == r_count_7_io_out ? io_r_104_b : _GEN_3083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3085 = 9'h69 == r_count_7_io_out ? io_r_105_b : _GEN_3084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3086 = 9'h6a == r_count_7_io_out ? io_r_106_b : _GEN_3085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3087 = 9'h6b == r_count_7_io_out ? io_r_107_b : _GEN_3086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3088 = 9'h6c == r_count_7_io_out ? io_r_108_b : _GEN_3087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3089 = 9'h6d == r_count_7_io_out ? io_r_109_b : _GEN_3088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3090 = 9'h6e == r_count_7_io_out ? io_r_110_b : _GEN_3089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3091 = 9'h6f == r_count_7_io_out ? io_r_111_b : _GEN_3090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3092 = 9'h70 == r_count_7_io_out ? io_r_112_b : _GEN_3091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3093 = 9'h71 == r_count_7_io_out ? io_r_113_b : _GEN_3092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3094 = 9'h72 == r_count_7_io_out ? io_r_114_b : _GEN_3093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3095 = 9'h73 == r_count_7_io_out ? io_r_115_b : _GEN_3094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3096 = 9'h74 == r_count_7_io_out ? io_r_116_b : _GEN_3095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3097 = 9'h75 == r_count_7_io_out ? io_r_117_b : _GEN_3096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3098 = 9'h76 == r_count_7_io_out ? io_r_118_b : _GEN_3097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3099 = 9'h77 == r_count_7_io_out ? io_r_119_b : _GEN_3098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3100 = 9'h78 == r_count_7_io_out ? io_r_120_b : _GEN_3099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3101 = 9'h79 == r_count_7_io_out ? io_r_121_b : _GEN_3100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3102 = 9'h7a == r_count_7_io_out ? io_r_122_b : _GEN_3101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3103 = 9'h7b == r_count_7_io_out ? io_r_123_b : _GEN_3102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3104 = 9'h7c == r_count_7_io_out ? io_r_124_b : _GEN_3103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3105 = 9'h7d == r_count_7_io_out ? io_r_125_b : _GEN_3104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3106 = 9'h7e == r_count_7_io_out ? io_r_126_b : _GEN_3105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3107 = 9'h7f == r_count_7_io_out ? io_r_127_b : _GEN_3106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3108 = 9'h80 == r_count_7_io_out ? io_r_128_b : _GEN_3107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3109 = 9'h81 == r_count_7_io_out ? io_r_129_b : _GEN_3108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3110 = 9'h82 == r_count_7_io_out ? io_r_130_b : _GEN_3109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3111 = 9'h83 == r_count_7_io_out ? io_r_131_b : _GEN_3110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3112 = 9'h84 == r_count_7_io_out ? io_r_132_b : _GEN_3111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3113 = 9'h85 == r_count_7_io_out ? io_r_133_b : _GEN_3112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3114 = 9'h86 == r_count_7_io_out ? io_r_134_b : _GEN_3113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3115 = 9'h87 == r_count_7_io_out ? io_r_135_b : _GEN_3114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3116 = 9'h88 == r_count_7_io_out ? io_r_136_b : _GEN_3115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3117 = 9'h89 == r_count_7_io_out ? io_r_137_b : _GEN_3116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3118 = 9'h8a == r_count_7_io_out ? io_r_138_b : _GEN_3117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3119 = 9'h8b == r_count_7_io_out ? io_r_139_b : _GEN_3118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3120 = 9'h8c == r_count_7_io_out ? io_r_140_b : _GEN_3119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3121 = 9'h8d == r_count_7_io_out ? io_r_141_b : _GEN_3120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3122 = 9'h8e == r_count_7_io_out ? io_r_142_b : _GEN_3121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3123 = 9'h8f == r_count_7_io_out ? io_r_143_b : _GEN_3122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3124 = 9'h90 == r_count_7_io_out ? io_r_144_b : _GEN_3123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3125 = 9'h91 == r_count_7_io_out ? io_r_145_b : _GEN_3124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3126 = 9'h92 == r_count_7_io_out ? io_r_146_b : _GEN_3125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3127 = 9'h93 == r_count_7_io_out ? io_r_147_b : _GEN_3126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3128 = 9'h94 == r_count_7_io_out ? io_r_148_b : _GEN_3127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3129 = 9'h95 == r_count_7_io_out ? io_r_149_b : _GEN_3128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3130 = 9'h96 == r_count_7_io_out ? io_r_150_b : _GEN_3129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3131 = 9'h97 == r_count_7_io_out ? io_r_151_b : _GEN_3130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3132 = 9'h98 == r_count_7_io_out ? io_r_152_b : _GEN_3131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3133 = 9'h99 == r_count_7_io_out ? io_r_153_b : _GEN_3132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3134 = 9'h9a == r_count_7_io_out ? io_r_154_b : _GEN_3133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3135 = 9'h9b == r_count_7_io_out ? io_r_155_b : _GEN_3134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3136 = 9'h9c == r_count_7_io_out ? io_r_156_b : _GEN_3135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3137 = 9'h9d == r_count_7_io_out ? io_r_157_b : _GEN_3136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3138 = 9'h9e == r_count_7_io_out ? io_r_158_b : _GEN_3137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3139 = 9'h9f == r_count_7_io_out ? io_r_159_b : _GEN_3138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3140 = 9'ha0 == r_count_7_io_out ? io_r_160_b : _GEN_3139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3141 = 9'ha1 == r_count_7_io_out ? io_r_161_b : _GEN_3140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3142 = 9'ha2 == r_count_7_io_out ? io_r_162_b : _GEN_3141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3143 = 9'ha3 == r_count_7_io_out ? io_r_163_b : _GEN_3142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3144 = 9'ha4 == r_count_7_io_out ? io_r_164_b : _GEN_3143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3145 = 9'ha5 == r_count_7_io_out ? io_r_165_b : _GEN_3144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3146 = 9'ha6 == r_count_7_io_out ? io_r_166_b : _GEN_3145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3147 = 9'ha7 == r_count_7_io_out ? io_r_167_b : _GEN_3146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3148 = 9'ha8 == r_count_7_io_out ? io_r_168_b : _GEN_3147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3149 = 9'ha9 == r_count_7_io_out ? io_r_169_b : _GEN_3148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3150 = 9'haa == r_count_7_io_out ? io_r_170_b : _GEN_3149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3151 = 9'hab == r_count_7_io_out ? io_r_171_b : _GEN_3150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3152 = 9'hac == r_count_7_io_out ? io_r_172_b : _GEN_3151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3153 = 9'had == r_count_7_io_out ? io_r_173_b : _GEN_3152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3154 = 9'hae == r_count_7_io_out ? io_r_174_b : _GEN_3153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3155 = 9'haf == r_count_7_io_out ? io_r_175_b : _GEN_3154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3156 = 9'hb0 == r_count_7_io_out ? io_r_176_b : _GEN_3155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3157 = 9'hb1 == r_count_7_io_out ? io_r_177_b : _GEN_3156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3158 = 9'hb2 == r_count_7_io_out ? io_r_178_b : _GEN_3157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3159 = 9'hb3 == r_count_7_io_out ? io_r_179_b : _GEN_3158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3160 = 9'hb4 == r_count_7_io_out ? io_r_180_b : _GEN_3159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3161 = 9'hb5 == r_count_7_io_out ? io_r_181_b : _GEN_3160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3162 = 9'hb6 == r_count_7_io_out ? io_r_182_b : _GEN_3161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3163 = 9'hb7 == r_count_7_io_out ? io_r_183_b : _GEN_3162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3164 = 9'hb8 == r_count_7_io_out ? io_r_184_b : _GEN_3163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3165 = 9'hb9 == r_count_7_io_out ? io_r_185_b : _GEN_3164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3166 = 9'hba == r_count_7_io_out ? io_r_186_b : _GEN_3165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3167 = 9'hbb == r_count_7_io_out ? io_r_187_b : _GEN_3166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3168 = 9'hbc == r_count_7_io_out ? io_r_188_b : _GEN_3167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3169 = 9'hbd == r_count_7_io_out ? io_r_189_b : _GEN_3168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3170 = 9'hbe == r_count_7_io_out ? io_r_190_b : _GEN_3169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3171 = 9'hbf == r_count_7_io_out ? io_r_191_b : _GEN_3170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3172 = 9'hc0 == r_count_7_io_out ? io_r_192_b : _GEN_3171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3173 = 9'hc1 == r_count_7_io_out ? io_r_193_b : _GEN_3172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3174 = 9'hc2 == r_count_7_io_out ? io_r_194_b : _GEN_3173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3175 = 9'hc3 == r_count_7_io_out ? io_r_195_b : _GEN_3174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3176 = 9'hc4 == r_count_7_io_out ? io_r_196_b : _GEN_3175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3177 = 9'hc5 == r_count_7_io_out ? io_r_197_b : _GEN_3176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3178 = 9'hc6 == r_count_7_io_out ? io_r_198_b : _GEN_3177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3179 = 9'hc7 == r_count_7_io_out ? io_r_199_b : _GEN_3178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3180 = 9'hc8 == r_count_7_io_out ? io_r_200_b : _GEN_3179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3181 = 9'hc9 == r_count_7_io_out ? io_r_201_b : _GEN_3180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3182 = 9'hca == r_count_7_io_out ? io_r_202_b : _GEN_3181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3183 = 9'hcb == r_count_7_io_out ? io_r_203_b : _GEN_3182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3184 = 9'hcc == r_count_7_io_out ? io_r_204_b : _GEN_3183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3185 = 9'hcd == r_count_7_io_out ? io_r_205_b : _GEN_3184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3186 = 9'hce == r_count_7_io_out ? io_r_206_b : _GEN_3185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3187 = 9'hcf == r_count_7_io_out ? io_r_207_b : _GEN_3186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3188 = 9'hd0 == r_count_7_io_out ? io_r_208_b : _GEN_3187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3189 = 9'hd1 == r_count_7_io_out ? io_r_209_b : _GEN_3188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3190 = 9'hd2 == r_count_7_io_out ? io_r_210_b : _GEN_3189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3191 = 9'hd3 == r_count_7_io_out ? io_r_211_b : _GEN_3190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3192 = 9'hd4 == r_count_7_io_out ? io_r_212_b : _GEN_3191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3193 = 9'hd5 == r_count_7_io_out ? io_r_213_b : _GEN_3192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3194 = 9'hd6 == r_count_7_io_out ? io_r_214_b : _GEN_3193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3195 = 9'hd7 == r_count_7_io_out ? io_r_215_b : _GEN_3194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3196 = 9'hd8 == r_count_7_io_out ? io_r_216_b : _GEN_3195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3197 = 9'hd9 == r_count_7_io_out ? io_r_217_b : _GEN_3196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3198 = 9'hda == r_count_7_io_out ? io_r_218_b : _GEN_3197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3199 = 9'hdb == r_count_7_io_out ? io_r_219_b : _GEN_3198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3200 = 9'hdc == r_count_7_io_out ? io_r_220_b : _GEN_3199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3201 = 9'hdd == r_count_7_io_out ? io_r_221_b : _GEN_3200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3202 = 9'hde == r_count_7_io_out ? io_r_222_b : _GEN_3201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3203 = 9'hdf == r_count_7_io_out ? io_r_223_b : _GEN_3202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3204 = 9'he0 == r_count_7_io_out ? io_r_224_b : _GEN_3203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3205 = 9'he1 == r_count_7_io_out ? io_r_225_b : _GEN_3204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3206 = 9'he2 == r_count_7_io_out ? io_r_226_b : _GEN_3205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3207 = 9'he3 == r_count_7_io_out ? io_r_227_b : _GEN_3206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3208 = 9'he4 == r_count_7_io_out ? io_r_228_b : _GEN_3207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3209 = 9'he5 == r_count_7_io_out ? io_r_229_b : _GEN_3208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3210 = 9'he6 == r_count_7_io_out ? io_r_230_b : _GEN_3209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3211 = 9'he7 == r_count_7_io_out ? io_r_231_b : _GEN_3210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3212 = 9'he8 == r_count_7_io_out ? io_r_232_b : _GEN_3211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3213 = 9'he9 == r_count_7_io_out ? io_r_233_b : _GEN_3212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3214 = 9'hea == r_count_7_io_out ? io_r_234_b : _GEN_3213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3215 = 9'heb == r_count_7_io_out ? io_r_235_b : _GEN_3214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3216 = 9'hec == r_count_7_io_out ? io_r_236_b : _GEN_3215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3217 = 9'hed == r_count_7_io_out ? io_r_237_b : _GEN_3216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3218 = 9'hee == r_count_7_io_out ? io_r_238_b : _GEN_3217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3219 = 9'hef == r_count_7_io_out ? io_r_239_b : _GEN_3218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3220 = 9'hf0 == r_count_7_io_out ? io_r_240_b : _GEN_3219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3221 = 9'hf1 == r_count_7_io_out ? io_r_241_b : _GEN_3220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3222 = 9'hf2 == r_count_7_io_out ? io_r_242_b : _GEN_3221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3223 = 9'hf3 == r_count_7_io_out ? io_r_243_b : _GEN_3222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3224 = 9'hf4 == r_count_7_io_out ? io_r_244_b : _GEN_3223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3225 = 9'hf5 == r_count_7_io_out ? io_r_245_b : _GEN_3224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3226 = 9'hf6 == r_count_7_io_out ? io_r_246_b : _GEN_3225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3227 = 9'hf7 == r_count_7_io_out ? io_r_247_b : _GEN_3226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3228 = 9'hf8 == r_count_7_io_out ? io_r_248_b : _GEN_3227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3229 = 9'hf9 == r_count_7_io_out ? io_r_249_b : _GEN_3228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3230 = 9'hfa == r_count_7_io_out ? io_r_250_b : _GEN_3229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3231 = 9'hfb == r_count_7_io_out ? io_r_251_b : _GEN_3230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3232 = 9'hfc == r_count_7_io_out ? io_r_252_b : _GEN_3231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3233 = 9'hfd == r_count_7_io_out ? io_r_253_b : _GEN_3232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3234 = 9'hfe == r_count_7_io_out ? io_r_254_b : _GEN_3233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3235 = 9'hff == r_count_7_io_out ? io_r_255_b : _GEN_3234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3236 = 9'h100 == r_count_7_io_out ? io_r_256_b : _GEN_3235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3237 = 9'h101 == r_count_7_io_out ? io_r_257_b : _GEN_3236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3238 = 9'h102 == r_count_7_io_out ? io_r_258_b : _GEN_3237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3239 = 9'h103 == r_count_7_io_out ? io_r_259_b : _GEN_3238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3240 = 9'h104 == r_count_7_io_out ? io_r_260_b : _GEN_3239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3241 = 9'h105 == r_count_7_io_out ? io_r_261_b : _GEN_3240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3242 = 9'h106 == r_count_7_io_out ? io_r_262_b : _GEN_3241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3243 = 9'h107 == r_count_7_io_out ? io_r_263_b : _GEN_3242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3244 = 9'h108 == r_count_7_io_out ? io_r_264_b : _GEN_3243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3245 = 9'h109 == r_count_7_io_out ? io_r_265_b : _GEN_3244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3246 = 9'h10a == r_count_7_io_out ? io_r_266_b : _GEN_3245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3247 = 9'h10b == r_count_7_io_out ? io_r_267_b : _GEN_3246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3248 = 9'h10c == r_count_7_io_out ? io_r_268_b : _GEN_3247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3249 = 9'h10d == r_count_7_io_out ? io_r_269_b : _GEN_3248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3250 = 9'h10e == r_count_7_io_out ? io_r_270_b : _GEN_3249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3251 = 9'h10f == r_count_7_io_out ? io_r_271_b : _GEN_3250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3252 = 9'h110 == r_count_7_io_out ? io_r_272_b : _GEN_3251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3253 = 9'h111 == r_count_7_io_out ? io_r_273_b : _GEN_3252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3254 = 9'h112 == r_count_7_io_out ? io_r_274_b : _GEN_3253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3255 = 9'h113 == r_count_7_io_out ? io_r_275_b : _GEN_3254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3256 = 9'h114 == r_count_7_io_out ? io_r_276_b : _GEN_3255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3257 = 9'h115 == r_count_7_io_out ? io_r_277_b : _GEN_3256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3258 = 9'h116 == r_count_7_io_out ? io_r_278_b : _GEN_3257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3259 = 9'h117 == r_count_7_io_out ? io_r_279_b : _GEN_3258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3260 = 9'h118 == r_count_7_io_out ? io_r_280_b : _GEN_3259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3261 = 9'h119 == r_count_7_io_out ? io_r_281_b : _GEN_3260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3262 = 9'h11a == r_count_7_io_out ? io_r_282_b : _GEN_3261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3263 = 9'h11b == r_count_7_io_out ? io_r_283_b : _GEN_3262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3264 = 9'h11c == r_count_7_io_out ? io_r_284_b : _GEN_3263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3265 = 9'h11d == r_count_7_io_out ? io_r_285_b : _GEN_3264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3266 = 9'h11e == r_count_7_io_out ? io_r_286_b : _GEN_3265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3267 = 9'h11f == r_count_7_io_out ? io_r_287_b : _GEN_3266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3268 = 9'h120 == r_count_7_io_out ? io_r_288_b : _GEN_3267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3269 = 9'h121 == r_count_7_io_out ? io_r_289_b : _GEN_3268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3270 = 9'h122 == r_count_7_io_out ? io_r_290_b : _GEN_3269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3271 = 9'h123 == r_count_7_io_out ? io_r_291_b : _GEN_3270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3272 = 9'h124 == r_count_7_io_out ? io_r_292_b : _GEN_3271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3273 = 9'h125 == r_count_7_io_out ? io_r_293_b : _GEN_3272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3274 = 9'h126 == r_count_7_io_out ? io_r_294_b : _GEN_3273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3275 = 9'h127 == r_count_7_io_out ? io_r_295_b : _GEN_3274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3276 = 9'h128 == r_count_7_io_out ? io_r_296_b : _GEN_3275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3277 = 9'h129 == r_count_7_io_out ? io_r_297_b : _GEN_3276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3278 = 9'h12a == r_count_7_io_out ? io_r_298_b : _GEN_3277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3279 = 9'h12b == r_count_7_io_out ? io_r_299_b : _GEN_3278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3280 = 9'h12c == r_count_7_io_out ? io_r_300_b : _GEN_3279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3281 = 9'h12d == r_count_7_io_out ? io_r_301_b : _GEN_3280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3282 = 9'h12e == r_count_7_io_out ? io_r_302_b : _GEN_3281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3283 = 9'h12f == r_count_7_io_out ? io_r_303_b : _GEN_3282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3284 = 9'h130 == r_count_7_io_out ? io_r_304_b : _GEN_3283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3285 = 9'h131 == r_count_7_io_out ? io_r_305_b : _GEN_3284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3286 = 9'h132 == r_count_7_io_out ? io_r_306_b : _GEN_3285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3287 = 9'h133 == r_count_7_io_out ? io_r_307_b : _GEN_3286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3288 = 9'h134 == r_count_7_io_out ? io_r_308_b : _GEN_3287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3289 = 9'h135 == r_count_7_io_out ? io_r_309_b : _GEN_3288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3290 = 9'h136 == r_count_7_io_out ? io_r_310_b : _GEN_3289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3291 = 9'h137 == r_count_7_io_out ? io_r_311_b : _GEN_3290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3292 = 9'h138 == r_count_7_io_out ? io_r_312_b : _GEN_3291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3293 = 9'h139 == r_count_7_io_out ? io_r_313_b : _GEN_3292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3294 = 9'h13a == r_count_7_io_out ? io_r_314_b : _GEN_3293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3295 = 9'h13b == r_count_7_io_out ? io_r_315_b : _GEN_3294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3296 = 9'h13c == r_count_7_io_out ? io_r_316_b : _GEN_3295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3297 = 9'h13d == r_count_7_io_out ? io_r_317_b : _GEN_3296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3298 = 9'h13e == r_count_7_io_out ? io_r_318_b : _GEN_3297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3299 = 9'h13f == r_count_7_io_out ? io_r_319_b : _GEN_3298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3300 = 9'h140 == r_count_7_io_out ? io_r_320_b : _GEN_3299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3301 = 9'h141 == r_count_7_io_out ? io_r_321_b : _GEN_3300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3302 = 9'h142 == r_count_7_io_out ? io_r_322_b : _GEN_3301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3303 = 9'h143 == r_count_7_io_out ? io_r_323_b : _GEN_3302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3304 = 9'h144 == r_count_7_io_out ? io_r_324_b : _GEN_3303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3305 = 9'h145 == r_count_7_io_out ? io_r_325_b : _GEN_3304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3306 = 9'h146 == r_count_7_io_out ? io_r_326_b : _GEN_3305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3307 = 9'h147 == r_count_7_io_out ? io_r_327_b : _GEN_3306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3308 = 9'h148 == r_count_7_io_out ? io_r_328_b : _GEN_3307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3309 = 9'h149 == r_count_7_io_out ? io_r_329_b : _GEN_3308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3310 = 9'h14a == r_count_7_io_out ? io_r_330_b : _GEN_3309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3311 = 9'h14b == r_count_7_io_out ? io_r_331_b : _GEN_3310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3312 = 9'h14c == r_count_7_io_out ? io_r_332_b : _GEN_3311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3313 = 9'h14d == r_count_7_io_out ? io_r_333_b : _GEN_3312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3314 = 9'h14e == r_count_7_io_out ? io_r_334_b : _GEN_3313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3315 = 9'h14f == r_count_7_io_out ? io_r_335_b : _GEN_3314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3316 = 9'h150 == r_count_7_io_out ? io_r_336_b : _GEN_3315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3317 = 9'h151 == r_count_7_io_out ? io_r_337_b : _GEN_3316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3318 = 9'h152 == r_count_7_io_out ? io_r_338_b : _GEN_3317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3319 = 9'h153 == r_count_7_io_out ? io_r_339_b : _GEN_3318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3320 = 9'h154 == r_count_7_io_out ? io_r_340_b : _GEN_3319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3321 = 9'h155 == r_count_7_io_out ? io_r_341_b : _GEN_3320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3322 = 9'h156 == r_count_7_io_out ? io_r_342_b : _GEN_3321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3323 = 9'h157 == r_count_7_io_out ? io_r_343_b : _GEN_3322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3324 = 9'h158 == r_count_7_io_out ? io_r_344_b : _GEN_3323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3325 = 9'h159 == r_count_7_io_out ? io_r_345_b : _GEN_3324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3326 = 9'h15a == r_count_7_io_out ? io_r_346_b : _GEN_3325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3327 = 9'h15b == r_count_7_io_out ? io_r_347_b : _GEN_3326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3328 = 9'h15c == r_count_7_io_out ? io_r_348_b : _GEN_3327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3329 = 9'h15d == r_count_7_io_out ? io_r_349_b : _GEN_3328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3330 = 9'h15e == r_count_7_io_out ? io_r_350_b : _GEN_3329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3331 = 9'h15f == r_count_7_io_out ? io_r_351_b : _GEN_3330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3332 = 9'h160 == r_count_7_io_out ? io_r_352_b : _GEN_3331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3333 = 9'h161 == r_count_7_io_out ? io_r_353_b : _GEN_3332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3334 = 9'h162 == r_count_7_io_out ? io_r_354_b : _GEN_3333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3335 = 9'h163 == r_count_7_io_out ? io_r_355_b : _GEN_3334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3336 = 9'h164 == r_count_7_io_out ? io_r_356_b : _GEN_3335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3337 = 9'h165 == r_count_7_io_out ? io_r_357_b : _GEN_3336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3338 = 9'h166 == r_count_7_io_out ? io_r_358_b : _GEN_3337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3339 = 9'h167 == r_count_7_io_out ? io_r_359_b : _GEN_3338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3340 = 9'h168 == r_count_7_io_out ? io_r_360_b : _GEN_3339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3341 = 9'h169 == r_count_7_io_out ? io_r_361_b : _GEN_3340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3342 = 9'h16a == r_count_7_io_out ? io_r_362_b : _GEN_3341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3343 = 9'h16b == r_count_7_io_out ? io_r_363_b : _GEN_3342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3344 = 9'h16c == r_count_7_io_out ? io_r_364_b : _GEN_3343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3345 = 9'h16d == r_count_7_io_out ? io_r_365_b : _GEN_3344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3346 = 9'h16e == r_count_7_io_out ? io_r_366_b : _GEN_3345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3347 = 9'h16f == r_count_7_io_out ? io_r_367_b : _GEN_3346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3348 = 9'h170 == r_count_7_io_out ? io_r_368_b : _GEN_3347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3349 = 9'h171 == r_count_7_io_out ? io_r_369_b : _GEN_3348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3350 = 9'h172 == r_count_7_io_out ? io_r_370_b : _GEN_3349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3351 = 9'h173 == r_count_7_io_out ? io_r_371_b : _GEN_3350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3352 = 9'h174 == r_count_7_io_out ? io_r_372_b : _GEN_3351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3353 = 9'h175 == r_count_7_io_out ? io_r_373_b : _GEN_3352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3354 = 9'h176 == r_count_7_io_out ? io_r_374_b : _GEN_3353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3355 = 9'h177 == r_count_7_io_out ? io_r_375_b : _GEN_3354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3356 = 9'h178 == r_count_7_io_out ? io_r_376_b : _GEN_3355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3357 = 9'h179 == r_count_7_io_out ? io_r_377_b : _GEN_3356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3358 = 9'h17a == r_count_7_io_out ? io_r_378_b : _GEN_3357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3359 = 9'h17b == r_count_7_io_out ? io_r_379_b : _GEN_3358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3360 = 9'h17c == r_count_7_io_out ? io_r_380_b : _GEN_3359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3361 = 9'h17d == r_count_7_io_out ? io_r_381_b : _GEN_3360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3362 = 9'h17e == r_count_7_io_out ? io_r_382_b : _GEN_3361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3363 = 9'h17f == r_count_7_io_out ? io_r_383_b : _GEN_3362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3364 = 9'h180 == r_count_7_io_out ? io_r_384_b : _GEN_3363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3365 = 9'h181 == r_count_7_io_out ? io_r_385_b : _GEN_3364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3366 = 9'h182 == r_count_7_io_out ? io_r_386_b : _GEN_3365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3367 = 9'h183 == r_count_7_io_out ? io_r_387_b : _GEN_3366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3368 = 9'h184 == r_count_7_io_out ? io_r_388_b : _GEN_3367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3369 = 9'h185 == r_count_7_io_out ? io_r_389_b : _GEN_3368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3370 = 9'h186 == r_count_7_io_out ? io_r_390_b : _GEN_3369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3371 = 9'h187 == r_count_7_io_out ? io_r_391_b : _GEN_3370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3372 = 9'h188 == r_count_7_io_out ? io_r_392_b : _GEN_3371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3373 = 9'h189 == r_count_7_io_out ? io_r_393_b : _GEN_3372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3374 = 9'h18a == r_count_7_io_out ? io_r_394_b : _GEN_3373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3375 = 9'h18b == r_count_7_io_out ? io_r_395_b : _GEN_3374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3376 = 9'h18c == r_count_7_io_out ? io_r_396_b : _GEN_3375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3377 = 9'h18d == r_count_7_io_out ? io_r_397_b : _GEN_3376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3378 = 9'h18e == r_count_7_io_out ? io_r_398_b : _GEN_3377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3381 = 9'h1 == r_count_8_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3382 = 9'h2 == r_count_8_io_out ? io_r_2_b : _GEN_3381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3383 = 9'h3 == r_count_8_io_out ? io_r_3_b : _GEN_3382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3384 = 9'h4 == r_count_8_io_out ? io_r_4_b : _GEN_3383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3385 = 9'h5 == r_count_8_io_out ? io_r_5_b : _GEN_3384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3386 = 9'h6 == r_count_8_io_out ? io_r_6_b : _GEN_3385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3387 = 9'h7 == r_count_8_io_out ? io_r_7_b : _GEN_3386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3388 = 9'h8 == r_count_8_io_out ? io_r_8_b : _GEN_3387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3389 = 9'h9 == r_count_8_io_out ? io_r_9_b : _GEN_3388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3390 = 9'ha == r_count_8_io_out ? io_r_10_b : _GEN_3389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3391 = 9'hb == r_count_8_io_out ? io_r_11_b : _GEN_3390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3392 = 9'hc == r_count_8_io_out ? io_r_12_b : _GEN_3391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3393 = 9'hd == r_count_8_io_out ? io_r_13_b : _GEN_3392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3394 = 9'he == r_count_8_io_out ? io_r_14_b : _GEN_3393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3395 = 9'hf == r_count_8_io_out ? io_r_15_b : _GEN_3394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3396 = 9'h10 == r_count_8_io_out ? io_r_16_b : _GEN_3395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3397 = 9'h11 == r_count_8_io_out ? io_r_17_b : _GEN_3396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3398 = 9'h12 == r_count_8_io_out ? io_r_18_b : _GEN_3397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3399 = 9'h13 == r_count_8_io_out ? io_r_19_b : _GEN_3398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3400 = 9'h14 == r_count_8_io_out ? io_r_20_b : _GEN_3399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3401 = 9'h15 == r_count_8_io_out ? io_r_21_b : _GEN_3400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3402 = 9'h16 == r_count_8_io_out ? io_r_22_b : _GEN_3401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3403 = 9'h17 == r_count_8_io_out ? io_r_23_b : _GEN_3402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3404 = 9'h18 == r_count_8_io_out ? io_r_24_b : _GEN_3403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3405 = 9'h19 == r_count_8_io_out ? io_r_25_b : _GEN_3404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3406 = 9'h1a == r_count_8_io_out ? io_r_26_b : _GEN_3405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3407 = 9'h1b == r_count_8_io_out ? io_r_27_b : _GEN_3406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3408 = 9'h1c == r_count_8_io_out ? io_r_28_b : _GEN_3407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3409 = 9'h1d == r_count_8_io_out ? io_r_29_b : _GEN_3408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3410 = 9'h1e == r_count_8_io_out ? io_r_30_b : _GEN_3409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3411 = 9'h1f == r_count_8_io_out ? io_r_31_b : _GEN_3410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3412 = 9'h20 == r_count_8_io_out ? io_r_32_b : _GEN_3411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3413 = 9'h21 == r_count_8_io_out ? io_r_33_b : _GEN_3412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3414 = 9'h22 == r_count_8_io_out ? io_r_34_b : _GEN_3413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3415 = 9'h23 == r_count_8_io_out ? io_r_35_b : _GEN_3414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3416 = 9'h24 == r_count_8_io_out ? io_r_36_b : _GEN_3415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3417 = 9'h25 == r_count_8_io_out ? io_r_37_b : _GEN_3416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3418 = 9'h26 == r_count_8_io_out ? io_r_38_b : _GEN_3417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3419 = 9'h27 == r_count_8_io_out ? io_r_39_b : _GEN_3418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3420 = 9'h28 == r_count_8_io_out ? io_r_40_b : _GEN_3419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3421 = 9'h29 == r_count_8_io_out ? io_r_41_b : _GEN_3420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3422 = 9'h2a == r_count_8_io_out ? io_r_42_b : _GEN_3421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3423 = 9'h2b == r_count_8_io_out ? io_r_43_b : _GEN_3422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3424 = 9'h2c == r_count_8_io_out ? io_r_44_b : _GEN_3423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3425 = 9'h2d == r_count_8_io_out ? io_r_45_b : _GEN_3424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3426 = 9'h2e == r_count_8_io_out ? io_r_46_b : _GEN_3425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3427 = 9'h2f == r_count_8_io_out ? io_r_47_b : _GEN_3426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3428 = 9'h30 == r_count_8_io_out ? io_r_48_b : _GEN_3427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3429 = 9'h31 == r_count_8_io_out ? io_r_49_b : _GEN_3428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3430 = 9'h32 == r_count_8_io_out ? io_r_50_b : _GEN_3429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3431 = 9'h33 == r_count_8_io_out ? io_r_51_b : _GEN_3430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3432 = 9'h34 == r_count_8_io_out ? io_r_52_b : _GEN_3431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3433 = 9'h35 == r_count_8_io_out ? io_r_53_b : _GEN_3432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3434 = 9'h36 == r_count_8_io_out ? io_r_54_b : _GEN_3433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3435 = 9'h37 == r_count_8_io_out ? io_r_55_b : _GEN_3434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3436 = 9'h38 == r_count_8_io_out ? io_r_56_b : _GEN_3435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3437 = 9'h39 == r_count_8_io_out ? io_r_57_b : _GEN_3436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3438 = 9'h3a == r_count_8_io_out ? io_r_58_b : _GEN_3437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3439 = 9'h3b == r_count_8_io_out ? io_r_59_b : _GEN_3438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3440 = 9'h3c == r_count_8_io_out ? io_r_60_b : _GEN_3439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3441 = 9'h3d == r_count_8_io_out ? io_r_61_b : _GEN_3440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3442 = 9'h3e == r_count_8_io_out ? io_r_62_b : _GEN_3441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3443 = 9'h3f == r_count_8_io_out ? io_r_63_b : _GEN_3442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3444 = 9'h40 == r_count_8_io_out ? io_r_64_b : _GEN_3443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3445 = 9'h41 == r_count_8_io_out ? io_r_65_b : _GEN_3444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3446 = 9'h42 == r_count_8_io_out ? io_r_66_b : _GEN_3445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3447 = 9'h43 == r_count_8_io_out ? io_r_67_b : _GEN_3446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3448 = 9'h44 == r_count_8_io_out ? io_r_68_b : _GEN_3447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3449 = 9'h45 == r_count_8_io_out ? io_r_69_b : _GEN_3448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3450 = 9'h46 == r_count_8_io_out ? io_r_70_b : _GEN_3449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3451 = 9'h47 == r_count_8_io_out ? io_r_71_b : _GEN_3450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3452 = 9'h48 == r_count_8_io_out ? io_r_72_b : _GEN_3451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3453 = 9'h49 == r_count_8_io_out ? io_r_73_b : _GEN_3452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3454 = 9'h4a == r_count_8_io_out ? io_r_74_b : _GEN_3453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3455 = 9'h4b == r_count_8_io_out ? io_r_75_b : _GEN_3454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3456 = 9'h4c == r_count_8_io_out ? io_r_76_b : _GEN_3455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3457 = 9'h4d == r_count_8_io_out ? io_r_77_b : _GEN_3456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3458 = 9'h4e == r_count_8_io_out ? io_r_78_b : _GEN_3457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3459 = 9'h4f == r_count_8_io_out ? io_r_79_b : _GEN_3458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3460 = 9'h50 == r_count_8_io_out ? io_r_80_b : _GEN_3459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3461 = 9'h51 == r_count_8_io_out ? io_r_81_b : _GEN_3460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3462 = 9'h52 == r_count_8_io_out ? io_r_82_b : _GEN_3461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3463 = 9'h53 == r_count_8_io_out ? io_r_83_b : _GEN_3462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3464 = 9'h54 == r_count_8_io_out ? io_r_84_b : _GEN_3463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3465 = 9'h55 == r_count_8_io_out ? io_r_85_b : _GEN_3464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3466 = 9'h56 == r_count_8_io_out ? io_r_86_b : _GEN_3465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3467 = 9'h57 == r_count_8_io_out ? io_r_87_b : _GEN_3466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3468 = 9'h58 == r_count_8_io_out ? io_r_88_b : _GEN_3467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3469 = 9'h59 == r_count_8_io_out ? io_r_89_b : _GEN_3468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3470 = 9'h5a == r_count_8_io_out ? io_r_90_b : _GEN_3469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3471 = 9'h5b == r_count_8_io_out ? io_r_91_b : _GEN_3470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3472 = 9'h5c == r_count_8_io_out ? io_r_92_b : _GEN_3471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3473 = 9'h5d == r_count_8_io_out ? io_r_93_b : _GEN_3472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3474 = 9'h5e == r_count_8_io_out ? io_r_94_b : _GEN_3473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3475 = 9'h5f == r_count_8_io_out ? io_r_95_b : _GEN_3474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3476 = 9'h60 == r_count_8_io_out ? io_r_96_b : _GEN_3475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3477 = 9'h61 == r_count_8_io_out ? io_r_97_b : _GEN_3476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3478 = 9'h62 == r_count_8_io_out ? io_r_98_b : _GEN_3477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3479 = 9'h63 == r_count_8_io_out ? io_r_99_b : _GEN_3478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3480 = 9'h64 == r_count_8_io_out ? io_r_100_b : _GEN_3479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3481 = 9'h65 == r_count_8_io_out ? io_r_101_b : _GEN_3480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3482 = 9'h66 == r_count_8_io_out ? io_r_102_b : _GEN_3481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3483 = 9'h67 == r_count_8_io_out ? io_r_103_b : _GEN_3482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3484 = 9'h68 == r_count_8_io_out ? io_r_104_b : _GEN_3483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3485 = 9'h69 == r_count_8_io_out ? io_r_105_b : _GEN_3484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3486 = 9'h6a == r_count_8_io_out ? io_r_106_b : _GEN_3485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3487 = 9'h6b == r_count_8_io_out ? io_r_107_b : _GEN_3486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3488 = 9'h6c == r_count_8_io_out ? io_r_108_b : _GEN_3487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3489 = 9'h6d == r_count_8_io_out ? io_r_109_b : _GEN_3488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3490 = 9'h6e == r_count_8_io_out ? io_r_110_b : _GEN_3489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3491 = 9'h6f == r_count_8_io_out ? io_r_111_b : _GEN_3490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3492 = 9'h70 == r_count_8_io_out ? io_r_112_b : _GEN_3491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3493 = 9'h71 == r_count_8_io_out ? io_r_113_b : _GEN_3492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3494 = 9'h72 == r_count_8_io_out ? io_r_114_b : _GEN_3493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3495 = 9'h73 == r_count_8_io_out ? io_r_115_b : _GEN_3494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3496 = 9'h74 == r_count_8_io_out ? io_r_116_b : _GEN_3495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3497 = 9'h75 == r_count_8_io_out ? io_r_117_b : _GEN_3496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3498 = 9'h76 == r_count_8_io_out ? io_r_118_b : _GEN_3497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3499 = 9'h77 == r_count_8_io_out ? io_r_119_b : _GEN_3498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3500 = 9'h78 == r_count_8_io_out ? io_r_120_b : _GEN_3499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3501 = 9'h79 == r_count_8_io_out ? io_r_121_b : _GEN_3500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3502 = 9'h7a == r_count_8_io_out ? io_r_122_b : _GEN_3501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3503 = 9'h7b == r_count_8_io_out ? io_r_123_b : _GEN_3502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3504 = 9'h7c == r_count_8_io_out ? io_r_124_b : _GEN_3503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3505 = 9'h7d == r_count_8_io_out ? io_r_125_b : _GEN_3504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3506 = 9'h7e == r_count_8_io_out ? io_r_126_b : _GEN_3505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3507 = 9'h7f == r_count_8_io_out ? io_r_127_b : _GEN_3506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3508 = 9'h80 == r_count_8_io_out ? io_r_128_b : _GEN_3507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3509 = 9'h81 == r_count_8_io_out ? io_r_129_b : _GEN_3508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3510 = 9'h82 == r_count_8_io_out ? io_r_130_b : _GEN_3509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3511 = 9'h83 == r_count_8_io_out ? io_r_131_b : _GEN_3510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3512 = 9'h84 == r_count_8_io_out ? io_r_132_b : _GEN_3511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3513 = 9'h85 == r_count_8_io_out ? io_r_133_b : _GEN_3512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3514 = 9'h86 == r_count_8_io_out ? io_r_134_b : _GEN_3513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3515 = 9'h87 == r_count_8_io_out ? io_r_135_b : _GEN_3514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3516 = 9'h88 == r_count_8_io_out ? io_r_136_b : _GEN_3515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3517 = 9'h89 == r_count_8_io_out ? io_r_137_b : _GEN_3516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3518 = 9'h8a == r_count_8_io_out ? io_r_138_b : _GEN_3517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3519 = 9'h8b == r_count_8_io_out ? io_r_139_b : _GEN_3518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3520 = 9'h8c == r_count_8_io_out ? io_r_140_b : _GEN_3519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3521 = 9'h8d == r_count_8_io_out ? io_r_141_b : _GEN_3520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3522 = 9'h8e == r_count_8_io_out ? io_r_142_b : _GEN_3521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3523 = 9'h8f == r_count_8_io_out ? io_r_143_b : _GEN_3522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3524 = 9'h90 == r_count_8_io_out ? io_r_144_b : _GEN_3523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3525 = 9'h91 == r_count_8_io_out ? io_r_145_b : _GEN_3524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3526 = 9'h92 == r_count_8_io_out ? io_r_146_b : _GEN_3525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3527 = 9'h93 == r_count_8_io_out ? io_r_147_b : _GEN_3526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3528 = 9'h94 == r_count_8_io_out ? io_r_148_b : _GEN_3527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3529 = 9'h95 == r_count_8_io_out ? io_r_149_b : _GEN_3528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3530 = 9'h96 == r_count_8_io_out ? io_r_150_b : _GEN_3529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3531 = 9'h97 == r_count_8_io_out ? io_r_151_b : _GEN_3530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3532 = 9'h98 == r_count_8_io_out ? io_r_152_b : _GEN_3531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3533 = 9'h99 == r_count_8_io_out ? io_r_153_b : _GEN_3532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3534 = 9'h9a == r_count_8_io_out ? io_r_154_b : _GEN_3533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3535 = 9'h9b == r_count_8_io_out ? io_r_155_b : _GEN_3534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3536 = 9'h9c == r_count_8_io_out ? io_r_156_b : _GEN_3535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3537 = 9'h9d == r_count_8_io_out ? io_r_157_b : _GEN_3536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3538 = 9'h9e == r_count_8_io_out ? io_r_158_b : _GEN_3537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3539 = 9'h9f == r_count_8_io_out ? io_r_159_b : _GEN_3538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3540 = 9'ha0 == r_count_8_io_out ? io_r_160_b : _GEN_3539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3541 = 9'ha1 == r_count_8_io_out ? io_r_161_b : _GEN_3540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3542 = 9'ha2 == r_count_8_io_out ? io_r_162_b : _GEN_3541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3543 = 9'ha3 == r_count_8_io_out ? io_r_163_b : _GEN_3542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3544 = 9'ha4 == r_count_8_io_out ? io_r_164_b : _GEN_3543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3545 = 9'ha5 == r_count_8_io_out ? io_r_165_b : _GEN_3544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3546 = 9'ha6 == r_count_8_io_out ? io_r_166_b : _GEN_3545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3547 = 9'ha7 == r_count_8_io_out ? io_r_167_b : _GEN_3546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3548 = 9'ha8 == r_count_8_io_out ? io_r_168_b : _GEN_3547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3549 = 9'ha9 == r_count_8_io_out ? io_r_169_b : _GEN_3548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3550 = 9'haa == r_count_8_io_out ? io_r_170_b : _GEN_3549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3551 = 9'hab == r_count_8_io_out ? io_r_171_b : _GEN_3550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3552 = 9'hac == r_count_8_io_out ? io_r_172_b : _GEN_3551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3553 = 9'had == r_count_8_io_out ? io_r_173_b : _GEN_3552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3554 = 9'hae == r_count_8_io_out ? io_r_174_b : _GEN_3553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3555 = 9'haf == r_count_8_io_out ? io_r_175_b : _GEN_3554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3556 = 9'hb0 == r_count_8_io_out ? io_r_176_b : _GEN_3555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3557 = 9'hb1 == r_count_8_io_out ? io_r_177_b : _GEN_3556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3558 = 9'hb2 == r_count_8_io_out ? io_r_178_b : _GEN_3557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3559 = 9'hb3 == r_count_8_io_out ? io_r_179_b : _GEN_3558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3560 = 9'hb4 == r_count_8_io_out ? io_r_180_b : _GEN_3559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3561 = 9'hb5 == r_count_8_io_out ? io_r_181_b : _GEN_3560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3562 = 9'hb6 == r_count_8_io_out ? io_r_182_b : _GEN_3561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3563 = 9'hb7 == r_count_8_io_out ? io_r_183_b : _GEN_3562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3564 = 9'hb8 == r_count_8_io_out ? io_r_184_b : _GEN_3563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3565 = 9'hb9 == r_count_8_io_out ? io_r_185_b : _GEN_3564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3566 = 9'hba == r_count_8_io_out ? io_r_186_b : _GEN_3565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3567 = 9'hbb == r_count_8_io_out ? io_r_187_b : _GEN_3566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3568 = 9'hbc == r_count_8_io_out ? io_r_188_b : _GEN_3567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3569 = 9'hbd == r_count_8_io_out ? io_r_189_b : _GEN_3568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3570 = 9'hbe == r_count_8_io_out ? io_r_190_b : _GEN_3569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3571 = 9'hbf == r_count_8_io_out ? io_r_191_b : _GEN_3570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3572 = 9'hc0 == r_count_8_io_out ? io_r_192_b : _GEN_3571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3573 = 9'hc1 == r_count_8_io_out ? io_r_193_b : _GEN_3572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3574 = 9'hc2 == r_count_8_io_out ? io_r_194_b : _GEN_3573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3575 = 9'hc3 == r_count_8_io_out ? io_r_195_b : _GEN_3574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3576 = 9'hc4 == r_count_8_io_out ? io_r_196_b : _GEN_3575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3577 = 9'hc5 == r_count_8_io_out ? io_r_197_b : _GEN_3576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3578 = 9'hc6 == r_count_8_io_out ? io_r_198_b : _GEN_3577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3579 = 9'hc7 == r_count_8_io_out ? io_r_199_b : _GEN_3578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3580 = 9'hc8 == r_count_8_io_out ? io_r_200_b : _GEN_3579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3581 = 9'hc9 == r_count_8_io_out ? io_r_201_b : _GEN_3580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3582 = 9'hca == r_count_8_io_out ? io_r_202_b : _GEN_3581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3583 = 9'hcb == r_count_8_io_out ? io_r_203_b : _GEN_3582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3584 = 9'hcc == r_count_8_io_out ? io_r_204_b : _GEN_3583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3585 = 9'hcd == r_count_8_io_out ? io_r_205_b : _GEN_3584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3586 = 9'hce == r_count_8_io_out ? io_r_206_b : _GEN_3585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3587 = 9'hcf == r_count_8_io_out ? io_r_207_b : _GEN_3586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3588 = 9'hd0 == r_count_8_io_out ? io_r_208_b : _GEN_3587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3589 = 9'hd1 == r_count_8_io_out ? io_r_209_b : _GEN_3588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3590 = 9'hd2 == r_count_8_io_out ? io_r_210_b : _GEN_3589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3591 = 9'hd3 == r_count_8_io_out ? io_r_211_b : _GEN_3590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3592 = 9'hd4 == r_count_8_io_out ? io_r_212_b : _GEN_3591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3593 = 9'hd5 == r_count_8_io_out ? io_r_213_b : _GEN_3592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3594 = 9'hd6 == r_count_8_io_out ? io_r_214_b : _GEN_3593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3595 = 9'hd7 == r_count_8_io_out ? io_r_215_b : _GEN_3594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3596 = 9'hd8 == r_count_8_io_out ? io_r_216_b : _GEN_3595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3597 = 9'hd9 == r_count_8_io_out ? io_r_217_b : _GEN_3596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3598 = 9'hda == r_count_8_io_out ? io_r_218_b : _GEN_3597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3599 = 9'hdb == r_count_8_io_out ? io_r_219_b : _GEN_3598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3600 = 9'hdc == r_count_8_io_out ? io_r_220_b : _GEN_3599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3601 = 9'hdd == r_count_8_io_out ? io_r_221_b : _GEN_3600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3602 = 9'hde == r_count_8_io_out ? io_r_222_b : _GEN_3601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3603 = 9'hdf == r_count_8_io_out ? io_r_223_b : _GEN_3602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3604 = 9'he0 == r_count_8_io_out ? io_r_224_b : _GEN_3603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3605 = 9'he1 == r_count_8_io_out ? io_r_225_b : _GEN_3604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3606 = 9'he2 == r_count_8_io_out ? io_r_226_b : _GEN_3605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3607 = 9'he3 == r_count_8_io_out ? io_r_227_b : _GEN_3606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3608 = 9'he4 == r_count_8_io_out ? io_r_228_b : _GEN_3607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3609 = 9'he5 == r_count_8_io_out ? io_r_229_b : _GEN_3608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3610 = 9'he6 == r_count_8_io_out ? io_r_230_b : _GEN_3609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3611 = 9'he7 == r_count_8_io_out ? io_r_231_b : _GEN_3610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3612 = 9'he8 == r_count_8_io_out ? io_r_232_b : _GEN_3611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3613 = 9'he9 == r_count_8_io_out ? io_r_233_b : _GEN_3612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3614 = 9'hea == r_count_8_io_out ? io_r_234_b : _GEN_3613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3615 = 9'heb == r_count_8_io_out ? io_r_235_b : _GEN_3614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3616 = 9'hec == r_count_8_io_out ? io_r_236_b : _GEN_3615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3617 = 9'hed == r_count_8_io_out ? io_r_237_b : _GEN_3616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3618 = 9'hee == r_count_8_io_out ? io_r_238_b : _GEN_3617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3619 = 9'hef == r_count_8_io_out ? io_r_239_b : _GEN_3618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3620 = 9'hf0 == r_count_8_io_out ? io_r_240_b : _GEN_3619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3621 = 9'hf1 == r_count_8_io_out ? io_r_241_b : _GEN_3620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3622 = 9'hf2 == r_count_8_io_out ? io_r_242_b : _GEN_3621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3623 = 9'hf3 == r_count_8_io_out ? io_r_243_b : _GEN_3622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3624 = 9'hf4 == r_count_8_io_out ? io_r_244_b : _GEN_3623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3625 = 9'hf5 == r_count_8_io_out ? io_r_245_b : _GEN_3624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3626 = 9'hf6 == r_count_8_io_out ? io_r_246_b : _GEN_3625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3627 = 9'hf7 == r_count_8_io_out ? io_r_247_b : _GEN_3626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3628 = 9'hf8 == r_count_8_io_out ? io_r_248_b : _GEN_3627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3629 = 9'hf9 == r_count_8_io_out ? io_r_249_b : _GEN_3628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3630 = 9'hfa == r_count_8_io_out ? io_r_250_b : _GEN_3629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3631 = 9'hfb == r_count_8_io_out ? io_r_251_b : _GEN_3630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3632 = 9'hfc == r_count_8_io_out ? io_r_252_b : _GEN_3631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3633 = 9'hfd == r_count_8_io_out ? io_r_253_b : _GEN_3632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3634 = 9'hfe == r_count_8_io_out ? io_r_254_b : _GEN_3633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3635 = 9'hff == r_count_8_io_out ? io_r_255_b : _GEN_3634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3636 = 9'h100 == r_count_8_io_out ? io_r_256_b : _GEN_3635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3637 = 9'h101 == r_count_8_io_out ? io_r_257_b : _GEN_3636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3638 = 9'h102 == r_count_8_io_out ? io_r_258_b : _GEN_3637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3639 = 9'h103 == r_count_8_io_out ? io_r_259_b : _GEN_3638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3640 = 9'h104 == r_count_8_io_out ? io_r_260_b : _GEN_3639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3641 = 9'h105 == r_count_8_io_out ? io_r_261_b : _GEN_3640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3642 = 9'h106 == r_count_8_io_out ? io_r_262_b : _GEN_3641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3643 = 9'h107 == r_count_8_io_out ? io_r_263_b : _GEN_3642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3644 = 9'h108 == r_count_8_io_out ? io_r_264_b : _GEN_3643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3645 = 9'h109 == r_count_8_io_out ? io_r_265_b : _GEN_3644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3646 = 9'h10a == r_count_8_io_out ? io_r_266_b : _GEN_3645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3647 = 9'h10b == r_count_8_io_out ? io_r_267_b : _GEN_3646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3648 = 9'h10c == r_count_8_io_out ? io_r_268_b : _GEN_3647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3649 = 9'h10d == r_count_8_io_out ? io_r_269_b : _GEN_3648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3650 = 9'h10e == r_count_8_io_out ? io_r_270_b : _GEN_3649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3651 = 9'h10f == r_count_8_io_out ? io_r_271_b : _GEN_3650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3652 = 9'h110 == r_count_8_io_out ? io_r_272_b : _GEN_3651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3653 = 9'h111 == r_count_8_io_out ? io_r_273_b : _GEN_3652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3654 = 9'h112 == r_count_8_io_out ? io_r_274_b : _GEN_3653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3655 = 9'h113 == r_count_8_io_out ? io_r_275_b : _GEN_3654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3656 = 9'h114 == r_count_8_io_out ? io_r_276_b : _GEN_3655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3657 = 9'h115 == r_count_8_io_out ? io_r_277_b : _GEN_3656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3658 = 9'h116 == r_count_8_io_out ? io_r_278_b : _GEN_3657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3659 = 9'h117 == r_count_8_io_out ? io_r_279_b : _GEN_3658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3660 = 9'h118 == r_count_8_io_out ? io_r_280_b : _GEN_3659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3661 = 9'h119 == r_count_8_io_out ? io_r_281_b : _GEN_3660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3662 = 9'h11a == r_count_8_io_out ? io_r_282_b : _GEN_3661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3663 = 9'h11b == r_count_8_io_out ? io_r_283_b : _GEN_3662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3664 = 9'h11c == r_count_8_io_out ? io_r_284_b : _GEN_3663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3665 = 9'h11d == r_count_8_io_out ? io_r_285_b : _GEN_3664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3666 = 9'h11e == r_count_8_io_out ? io_r_286_b : _GEN_3665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3667 = 9'h11f == r_count_8_io_out ? io_r_287_b : _GEN_3666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3668 = 9'h120 == r_count_8_io_out ? io_r_288_b : _GEN_3667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3669 = 9'h121 == r_count_8_io_out ? io_r_289_b : _GEN_3668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3670 = 9'h122 == r_count_8_io_out ? io_r_290_b : _GEN_3669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3671 = 9'h123 == r_count_8_io_out ? io_r_291_b : _GEN_3670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3672 = 9'h124 == r_count_8_io_out ? io_r_292_b : _GEN_3671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3673 = 9'h125 == r_count_8_io_out ? io_r_293_b : _GEN_3672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3674 = 9'h126 == r_count_8_io_out ? io_r_294_b : _GEN_3673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3675 = 9'h127 == r_count_8_io_out ? io_r_295_b : _GEN_3674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3676 = 9'h128 == r_count_8_io_out ? io_r_296_b : _GEN_3675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3677 = 9'h129 == r_count_8_io_out ? io_r_297_b : _GEN_3676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3678 = 9'h12a == r_count_8_io_out ? io_r_298_b : _GEN_3677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3679 = 9'h12b == r_count_8_io_out ? io_r_299_b : _GEN_3678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3680 = 9'h12c == r_count_8_io_out ? io_r_300_b : _GEN_3679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3681 = 9'h12d == r_count_8_io_out ? io_r_301_b : _GEN_3680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3682 = 9'h12e == r_count_8_io_out ? io_r_302_b : _GEN_3681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3683 = 9'h12f == r_count_8_io_out ? io_r_303_b : _GEN_3682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3684 = 9'h130 == r_count_8_io_out ? io_r_304_b : _GEN_3683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3685 = 9'h131 == r_count_8_io_out ? io_r_305_b : _GEN_3684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3686 = 9'h132 == r_count_8_io_out ? io_r_306_b : _GEN_3685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3687 = 9'h133 == r_count_8_io_out ? io_r_307_b : _GEN_3686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3688 = 9'h134 == r_count_8_io_out ? io_r_308_b : _GEN_3687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3689 = 9'h135 == r_count_8_io_out ? io_r_309_b : _GEN_3688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3690 = 9'h136 == r_count_8_io_out ? io_r_310_b : _GEN_3689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3691 = 9'h137 == r_count_8_io_out ? io_r_311_b : _GEN_3690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3692 = 9'h138 == r_count_8_io_out ? io_r_312_b : _GEN_3691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3693 = 9'h139 == r_count_8_io_out ? io_r_313_b : _GEN_3692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3694 = 9'h13a == r_count_8_io_out ? io_r_314_b : _GEN_3693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3695 = 9'h13b == r_count_8_io_out ? io_r_315_b : _GEN_3694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3696 = 9'h13c == r_count_8_io_out ? io_r_316_b : _GEN_3695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3697 = 9'h13d == r_count_8_io_out ? io_r_317_b : _GEN_3696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3698 = 9'h13e == r_count_8_io_out ? io_r_318_b : _GEN_3697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3699 = 9'h13f == r_count_8_io_out ? io_r_319_b : _GEN_3698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3700 = 9'h140 == r_count_8_io_out ? io_r_320_b : _GEN_3699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3701 = 9'h141 == r_count_8_io_out ? io_r_321_b : _GEN_3700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3702 = 9'h142 == r_count_8_io_out ? io_r_322_b : _GEN_3701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3703 = 9'h143 == r_count_8_io_out ? io_r_323_b : _GEN_3702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3704 = 9'h144 == r_count_8_io_out ? io_r_324_b : _GEN_3703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3705 = 9'h145 == r_count_8_io_out ? io_r_325_b : _GEN_3704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3706 = 9'h146 == r_count_8_io_out ? io_r_326_b : _GEN_3705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3707 = 9'h147 == r_count_8_io_out ? io_r_327_b : _GEN_3706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3708 = 9'h148 == r_count_8_io_out ? io_r_328_b : _GEN_3707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3709 = 9'h149 == r_count_8_io_out ? io_r_329_b : _GEN_3708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3710 = 9'h14a == r_count_8_io_out ? io_r_330_b : _GEN_3709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3711 = 9'h14b == r_count_8_io_out ? io_r_331_b : _GEN_3710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3712 = 9'h14c == r_count_8_io_out ? io_r_332_b : _GEN_3711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3713 = 9'h14d == r_count_8_io_out ? io_r_333_b : _GEN_3712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3714 = 9'h14e == r_count_8_io_out ? io_r_334_b : _GEN_3713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3715 = 9'h14f == r_count_8_io_out ? io_r_335_b : _GEN_3714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3716 = 9'h150 == r_count_8_io_out ? io_r_336_b : _GEN_3715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3717 = 9'h151 == r_count_8_io_out ? io_r_337_b : _GEN_3716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3718 = 9'h152 == r_count_8_io_out ? io_r_338_b : _GEN_3717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3719 = 9'h153 == r_count_8_io_out ? io_r_339_b : _GEN_3718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3720 = 9'h154 == r_count_8_io_out ? io_r_340_b : _GEN_3719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3721 = 9'h155 == r_count_8_io_out ? io_r_341_b : _GEN_3720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3722 = 9'h156 == r_count_8_io_out ? io_r_342_b : _GEN_3721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3723 = 9'h157 == r_count_8_io_out ? io_r_343_b : _GEN_3722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3724 = 9'h158 == r_count_8_io_out ? io_r_344_b : _GEN_3723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3725 = 9'h159 == r_count_8_io_out ? io_r_345_b : _GEN_3724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3726 = 9'h15a == r_count_8_io_out ? io_r_346_b : _GEN_3725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3727 = 9'h15b == r_count_8_io_out ? io_r_347_b : _GEN_3726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3728 = 9'h15c == r_count_8_io_out ? io_r_348_b : _GEN_3727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3729 = 9'h15d == r_count_8_io_out ? io_r_349_b : _GEN_3728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3730 = 9'h15e == r_count_8_io_out ? io_r_350_b : _GEN_3729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3731 = 9'h15f == r_count_8_io_out ? io_r_351_b : _GEN_3730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3732 = 9'h160 == r_count_8_io_out ? io_r_352_b : _GEN_3731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3733 = 9'h161 == r_count_8_io_out ? io_r_353_b : _GEN_3732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3734 = 9'h162 == r_count_8_io_out ? io_r_354_b : _GEN_3733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3735 = 9'h163 == r_count_8_io_out ? io_r_355_b : _GEN_3734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3736 = 9'h164 == r_count_8_io_out ? io_r_356_b : _GEN_3735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3737 = 9'h165 == r_count_8_io_out ? io_r_357_b : _GEN_3736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3738 = 9'h166 == r_count_8_io_out ? io_r_358_b : _GEN_3737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3739 = 9'h167 == r_count_8_io_out ? io_r_359_b : _GEN_3738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3740 = 9'h168 == r_count_8_io_out ? io_r_360_b : _GEN_3739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3741 = 9'h169 == r_count_8_io_out ? io_r_361_b : _GEN_3740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3742 = 9'h16a == r_count_8_io_out ? io_r_362_b : _GEN_3741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3743 = 9'h16b == r_count_8_io_out ? io_r_363_b : _GEN_3742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3744 = 9'h16c == r_count_8_io_out ? io_r_364_b : _GEN_3743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3745 = 9'h16d == r_count_8_io_out ? io_r_365_b : _GEN_3744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3746 = 9'h16e == r_count_8_io_out ? io_r_366_b : _GEN_3745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3747 = 9'h16f == r_count_8_io_out ? io_r_367_b : _GEN_3746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3748 = 9'h170 == r_count_8_io_out ? io_r_368_b : _GEN_3747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3749 = 9'h171 == r_count_8_io_out ? io_r_369_b : _GEN_3748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3750 = 9'h172 == r_count_8_io_out ? io_r_370_b : _GEN_3749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3751 = 9'h173 == r_count_8_io_out ? io_r_371_b : _GEN_3750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3752 = 9'h174 == r_count_8_io_out ? io_r_372_b : _GEN_3751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3753 = 9'h175 == r_count_8_io_out ? io_r_373_b : _GEN_3752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3754 = 9'h176 == r_count_8_io_out ? io_r_374_b : _GEN_3753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3755 = 9'h177 == r_count_8_io_out ? io_r_375_b : _GEN_3754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3756 = 9'h178 == r_count_8_io_out ? io_r_376_b : _GEN_3755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3757 = 9'h179 == r_count_8_io_out ? io_r_377_b : _GEN_3756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3758 = 9'h17a == r_count_8_io_out ? io_r_378_b : _GEN_3757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3759 = 9'h17b == r_count_8_io_out ? io_r_379_b : _GEN_3758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3760 = 9'h17c == r_count_8_io_out ? io_r_380_b : _GEN_3759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3761 = 9'h17d == r_count_8_io_out ? io_r_381_b : _GEN_3760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3762 = 9'h17e == r_count_8_io_out ? io_r_382_b : _GEN_3761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3763 = 9'h17f == r_count_8_io_out ? io_r_383_b : _GEN_3762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3764 = 9'h180 == r_count_8_io_out ? io_r_384_b : _GEN_3763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3765 = 9'h181 == r_count_8_io_out ? io_r_385_b : _GEN_3764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3766 = 9'h182 == r_count_8_io_out ? io_r_386_b : _GEN_3765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3767 = 9'h183 == r_count_8_io_out ? io_r_387_b : _GEN_3766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3768 = 9'h184 == r_count_8_io_out ? io_r_388_b : _GEN_3767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3769 = 9'h185 == r_count_8_io_out ? io_r_389_b : _GEN_3768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3770 = 9'h186 == r_count_8_io_out ? io_r_390_b : _GEN_3769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3771 = 9'h187 == r_count_8_io_out ? io_r_391_b : _GEN_3770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3772 = 9'h188 == r_count_8_io_out ? io_r_392_b : _GEN_3771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3773 = 9'h189 == r_count_8_io_out ? io_r_393_b : _GEN_3772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3774 = 9'h18a == r_count_8_io_out ? io_r_394_b : _GEN_3773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3775 = 9'h18b == r_count_8_io_out ? io_r_395_b : _GEN_3774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3776 = 9'h18c == r_count_8_io_out ? io_r_396_b : _GEN_3775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3777 = 9'h18d == r_count_8_io_out ? io_r_397_b : _GEN_3776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3778 = 9'h18e == r_count_8_io_out ? io_r_398_b : _GEN_3777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3781 = 9'h1 == r_count_9_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3782 = 9'h2 == r_count_9_io_out ? io_r_2_b : _GEN_3781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3783 = 9'h3 == r_count_9_io_out ? io_r_3_b : _GEN_3782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3784 = 9'h4 == r_count_9_io_out ? io_r_4_b : _GEN_3783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3785 = 9'h5 == r_count_9_io_out ? io_r_5_b : _GEN_3784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3786 = 9'h6 == r_count_9_io_out ? io_r_6_b : _GEN_3785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3787 = 9'h7 == r_count_9_io_out ? io_r_7_b : _GEN_3786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3788 = 9'h8 == r_count_9_io_out ? io_r_8_b : _GEN_3787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3789 = 9'h9 == r_count_9_io_out ? io_r_9_b : _GEN_3788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3790 = 9'ha == r_count_9_io_out ? io_r_10_b : _GEN_3789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3791 = 9'hb == r_count_9_io_out ? io_r_11_b : _GEN_3790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3792 = 9'hc == r_count_9_io_out ? io_r_12_b : _GEN_3791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3793 = 9'hd == r_count_9_io_out ? io_r_13_b : _GEN_3792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3794 = 9'he == r_count_9_io_out ? io_r_14_b : _GEN_3793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3795 = 9'hf == r_count_9_io_out ? io_r_15_b : _GEN_3794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3796 = 9'h10 == r_count_9_io_out ? io_r_16_b : _GEN_3795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3797 = 9'h11 == r_count_9_io_out ? io_r_17_b : _GEN_3796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3798 = 9'h12 == r_count_9_io_out ? io_r_18_b : _GEN_3797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3799 = 9'h13 == r_count_9_io_out ? io_r_19_b : _GEN_3798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3800 = 9'h14 == r_count_9_io_out ? io_r_20_b : _GEN_3799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3801 = 9'h15 == r_count_9_io_out ? io_r_21_b : _GEN_3800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3802 = 9'h16 == r_count_9_io_out ? io_r_22_b : _GEN_3801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3803 = 9'h17 == r_count_9_io_out ? io_r_23_b : _GEN_3802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3804 = 9'h18 == r_count_9_io_out ? io_r_24_b : _GEN_3803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3805 = 9'h19 == r_count_9_io_out ? io_r_25_b : _GEN_3804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3806 = 9'h1a == r_count_9_io_out ? io_r_26_b : _GEN_3805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3807 = 9'h1b == r_count_9_io_out ? io_r_27_b : _GEN_3806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3808 = 9'h1c == r_count_9_io_out ? io_r_28_b : _GEN_3807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3809 = 9'h1d == r_count_9_io_out ? io_r_29_b : _GEN_3808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3810 = 9'h1e == r_count_9_io_out ? io_r_30_b : _GEN_3809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3811 = 9'h1f == r_count_9_io_out ? io_r_31_b : _GEN_3810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3812 = 9'h20 == r_count_9_io_out ? io_r_32_b : _GEN_3811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3813 = 9'h21 == r_count_9_io_out ? io_r_33_b : _GEN_3812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3814 = 9'h22 == r_count_9_io_out ? io_r_34_b : _GEN_3813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3815 = 9'h23 == r_count_9_io_out ? io_r_35_b : _GEN_3814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3816 = 9'h24 == r_count_9_io_out ? io_r_36_b : _GEN_3815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3817 = 9'h25 == r_count_9_io_out ? io_r_37_b : _GEN_3816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3818 = 9'h26 == r_count_9_io_out ? io_r_38_b : _GEN_3817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3819 = 9'h27 == r_count_9_io_out ? io_r_39_b : _GEN_3818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3820 = 9'h28 == r_count_9_io_out ? io_r_40_b : _GEN_3819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3821 = 9'h29 == r_count_9_io_out ? io_r_41_b : _GEN_3820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3822 = 9'h2a == r_count_9_io_out ? io_r_42_b : _GEN_3821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3823 = 9'h2b == r_count_9_io_out ? io_r_43_b : _GEN_3822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3824 = 9'h2c == r_count_9_io_out ? io_r_44_b : _GEN_3823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3825 = 9'h2d == r_count_9_io_out ? io_r_45_b : _GEN_3824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3826 = 9'h2e == r_count_9_io_out ? io_r_46_b : _GEN_3825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3827 = 9'h2f == r_count_9_io_out ? io_r_47_b : _GEN_3826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3828 = 9'h30 == r_count_9_io_out ? io_r_48_b : _GEN_3827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3829 = 9'h31 == r_count_9_io_out ? io_r_49_b : _GEN_3828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3830 = 9'h32 == r_count_9_io_out ? io_r_50_b : _GEN_3829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3831 = 9'h33 == r_count_9_io_out ? io_r_51_b : _GEN_3830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3832 = 9'h34 == r_count_9_io_out ? io_r_52_b : _GEN_3831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3833 = 9'h35 == r_count_9_io_out ? io_r_53_b : _GEN_3832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3834 = 9'h36 == r_count_9_io_out ? io_r_54_b : _GEN_3833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3835 = 9'h37 == r_count_9_io_out ? io_r_55_b : _GEN_3834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3836 = 9'h38 == r_count_9_io_out ? io_r_56_b : _GEN_3835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3837 = 9'h39 == r_count_9_io_out ? io_r_57_b : _GEN_3836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3838 = 9'h3a == r_count_9_io_out ? io_r_58_b : _GEN_3837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3839 = 9'h3b == r_count_9_io_out ? io_r_59_b : _GEN_3838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3840 = 9'h3c == r_count_9_io_out ? io_r_60_b : _GEN_3839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3841 = 9'h3d == r_count_9_io_out ? io_r_61_b : _GEN_3840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3842 = 9'h3e == r_count_9_io_out ? io_r_62_b : _GEN_3841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3843 = 9'h3f == r_count_9_io_out ? io_r_63_b : _GEN_3842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3844 = 9'h40 == r_count_9_io_out ? io_r_64_b : _GEN_3843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3845 = 9'h41 == r_count_9_io_out ? io_r_65_b : _GEN_3844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3846 = 9'h42 == r_count_9_io_out ? io_r_66_b : _GEN_3845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3847 = 9'h43 == r_count_9_io_out ? io_r_67_b : _GEN_3846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3848 = 9'h44 == r_count_9_io_out ? io_r_68_b : _GEN_3847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3849 = 9'h45 == r_count_9_io_out ? io_r_69_b : _GEN_3848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3850 = 9'h46 == r_count_9_io_out ? io_r_70_b : _GEN_3849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3851 = 9'h47 == r_count_9_io_out ? io_r_71_b : _GEN_3850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3852 = 9'h48 == r_count_9_io_out ? io_r_72_b : _GEN_3851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3853 = 9'h49 == r_count_9_io_out ? io_r_73_b : _GEN_3852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3854 = 9'h4a == r_count_9_io_out ? io_r_74_b : _GEN_3853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3855 = 9'h4b == r_count_9_io_out ? io_r_75_b : _GEN_3854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3856 = 9'h4c == r_count_9_io_out ? io_r_76_b : _GEN_3855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3857 = 9'h4d == r_count_9_io_out ? io_r_77_b : _GEN_3856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3858 = 9'h4e == r_count_9_io_out ? io_r_78_b : _GEN_3857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3859 = 9'h4f == r_count_9_io_out ? io_r_79_b : _GEN_3858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3860 = 9'h50 == r_count_9_io_out ? io_r_80_b : _GEN_3859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3861 = 9'h51 == r_count_9_io_out ? io_r_81_b : _GEN_3860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3862 = 9'h52 == r_count_9_io_out ? io_r_82_b : _GEN_3861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3863 = 9'h53 == r_count_9_io_out ? io_r_83_b : _GEN_3862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3864 = 9'h54 == r_count_9_io_out ? io_r_84_b : _GEN_3863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3865 = 9'h55 == r_count_9_io_out ? io_r_85_b : _GEN_3864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3866 = 9'h56 == r_count_9_io_out ? io_r_86_b : _GEN_3865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3867 = 9'h57 == r_count_9_io_out ? io_r_87_b : _GEN_3866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3868 = 9'h58 == r_count_9_io_out ? io_r_88_b : _GEN_3867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3869 = 9'h59 == r_count_9_io_out ? io_r_89_b : _GEN_3868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3870 = 9'h5a == r_count_9_io_out ? io_r_90_b : _GEN_3869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3871 = 9'h5b == r_count_9_io_out ? io_r_91_b : _GEN_3870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3872 = 9'h5c == r_count_9_io_out ? io_r_92_b : _GEN_3871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3873 = 9'h5d == r_count_9_io_out ? io_r_93_b : _GEN_3872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3874 = 9'h5e == r_count_9_io_out ? io_r_94_b : _GEN_3873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3875 = 9'h5f == r_count_9_io_out ? io_r_95_b : _GEN_3874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3876 = 9'h60 == r_count_9_io_out ? io_r_96_b : _GEN_3875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3877 = 9'h61 == r_count_9_io_out ? io_r_97_b : _GEN_3876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3878 = 9'h62 == r_count_9_io_out ? io_r_98_b : _GEN_3877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3879 = 9'h63 == r_count_9_io_out ? io_r_99_b : _GEN_3878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3880 = 9'h64 == r_count_9_io_out ? io_r_100_b : _GEN_3879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3881 = 9'h65 == r_count_9_io_out ? io_r_101_b : _GEN_3880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3882 = 9'h66 == r_count_9_io_out ? io_r_102_b : _GEN_3881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3883 = 9'h67 == r_count_9_io_out ? io_r_103_b : _GEN_3882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3884 = 9'h68 == r_count_9_io_out ? io_r_104_b : _GEN_3883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3885 = 9'h69 == r_count_9_io_out ? io_r_105_b : _GEN_3884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3886 = 9'h6a == r_count_9_io_out ? io_r_106_b : _GEN_3885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3887 = 9'h6b == r_count_9_io_out ? io_r_107_b : _GEN_3886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3888 = 9'h6c == r_count_9_io_out ? io_r_108_b : _GEN_3887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3889 = 9'h6d == r_count_9_io_out ? io_r_109_b : _GEN_3888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3890 = 9'h6e == r_count_9_io_out ? io_r_110_b : _GEN_3889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3891 = 9'h6f == r_count_9_io_out ? io_r_111_b : _GEN_3890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3892 = 9'h70 == r_count_9_io_out ? io_r_112_b : _GEN_3891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3893 = 9'h71 == r_count_9_io_out ? io_r_113_b : _GEN_3892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3894 = 9'h72 == r_count_9_io_out ? io_r_114_b : _GEN_3893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3895 = 9'h73 == r_count_9_io_out ? io_r_115_b : _GEN_3894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3896 = 9'h74 == r_count_9_io_out ? io_r_116_b : _GEN_3895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3897 = 9'h75 == r_count_9_io_out ? io_r_117_b : _GEN_3896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3898 = 9'h76 == r_count_9_io_out ? io_r_118_b : _GEN_3897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3899 = 9'h77 == r_count_9_io_out ? io_r_119_b : _GEN_3898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3900 = 9'h78 == r_count_9_io_out ? io_r_120_b : _GEN_3899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3901 = 9'h79 == r_count_9_io_out ? io_r_121_b : _GEN_3900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3902 = 9'h7a == r_count_9_io_out ? io_r_122_b : _GEN_3901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3903 = 9'h7b == r_count_9_io_out ? io_r_123_b : _GEN_3902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3904 = 9'h7c == r_count_9_io_out ? io_r_124_b : _GEN_3903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3905 = 9'h7d == r_count_9_io_out ? io_r_125_b : _GEN_3904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3906 = 9'h7e == r_count_9_io_out ? io_r_126_b : _GEN_3905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3907 = 9'h7f == r_count_9_io_out ? io_r_127_b : _GEN_3906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3908 = 9'h80 == r_count_9_io_out ? io_r_128_b : _GEN_3907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3909 = 9'h81 == r_count_9_io_out ? io_r_129_b : _GEN_3908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3910 = 9'h82 == r_count_9_io_out ? io_r_130_b : _GEN_3909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3911 = 9'h83 == r_count_9_io_out ? io_r_131_b : _GEN_3910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3912 = 9'h84 == r_count_9_io_out ? io_r_132_b : _GEN_3911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3913 = 9'h85 == r_count_9_io_out ? io_r_133_b : _GEN_3912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3914 = 9'h86 == r_count_9_io_out ? io_r_134_b : _GEN_3913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3915 = 9'h87 == r_count_9_io_out ? io_r_135_b : _GEN_3914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3916 = 9'h88 == r_count_9_io_out ? io_r_136_b : _GEN_3915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3917 = 9'h89 == r_count_9_io_out ? io_r_137_b : _GEN_3916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3918 = 9'h8a == r_count_9_io_out ? io_r_138_b : _GEN_3917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3919 = 9'h8b == r_count_9_io_out ? io_r_139_b : _GEN_3918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3920 = 9'h8c == r_count_9_io_out ? io_r_140_b : _GEN_3919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3921 = 9'h8d == r_count_9_io_out ? io_r_141_b : _GEN_3920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3922 = 9'h8e == r_count_9_io_out ? io_r_142_b : _GEN_3921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3923 = 9'h8f == r_count_9_io_out ? io_r_143_b : _GEN_3922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3924 = 9'h90 == r_count_9_io_out ? io_r_144_b : _GEN_3923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3925 = 9'h91 == r_count_9_io_out ? io_r_145_b : _GEN_3924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3926 = 9'h92 == r_count_9_io_out ? io_r_146_b : _GEN_3925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3927 = 9'h93 == r_count_9_io_out ? io_r_147_b : _GEN_3926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3928 = 9'h94 == r_count_9_io_out ? io_r_148_b : _GEN_3927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3929 = 9'h95 == r_count_9_io_out ? io_r_149_b : _GEN_3928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3930 = 9'h96 == r_count_9_io_out ? io_r_150_b : _GEN_3929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3931 = 9'h97 == r_count_9_io_out ? io_r_151_b : _GEN_3930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3932 = 9'h98 == r_count_9_io_out ? io_r_152_b : _GEN_3931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3933 = 9'h99 == r_count_9_io_out ? io_r_153_b : _GEN_3932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3934 = 9'h9a == r_count_9_io_out ? io_r_154_b : _GEN_3933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3935 = 9'h9b == r_count_9_io_out ? io_r_155_b : _GEN_3934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3936 = 9'h9c == r_count_9_io_out ? io_r_156_b : _GEN_3935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3937 = 9'h9d == r_count_9_io_out ? io_r_157_b : _GEN_3936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3938 = 9'h9e == r_count_9_io_out ? io_r_158_b : _GEN_3937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3939 = 9'h9f == r_count_9_io_out ? io_r_159_b : _GEN_3938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3940 = 9'ha0 == r_count_9_io_out ? io_r_160_b : _GEN_3939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3941 = 9'ha1 == r_count_9_io_out ? io_r_161_b : _GEN_3940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3942 = 9'ha2 == r_count_9_io_out ? io_r_162_b : _GEN_3941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3943 = 9'ha3 == r_count_9_io_out ? io_r_163_b : _GEN_3942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3944 = 9'ha4 == r_count_9_io_out ? io_r_164_b : _GEN_3943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3945 = 9'ha5 == r_count_9_io_out ? io_r_165_b : _GEN_3944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3946 = 9'ha6 == r_count_9_io_out ? io_r_166_b : _GEN_3945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3947 = 9'ha7 == r_count_9_io_out ? io_r_167_b : _GEN_3946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3948 = 9'ha8 == r_count_9_io_out ? io_r_168_b : _GEN_3947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3949 = 9'ha9 == r_count_9_io_out ? io_r_169_b : _GEN_3948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3950 = 9'haa == r_count_9_io_out ? io_r_170_b : _GEN_3949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3951 = 9'hab == r_count_9_io_out ? io_r_171_b : _GEN_3950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3952 = 9'hac == r_count_9_io_out ? io_r_172_b : _GEN_3951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3953 = 9'had == r_count_9_io_out ? io_r_173_b : _GEN_3952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3954 = 9'hae == r_count_9_io_out ? io_r_174_b : _GEN_3953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3955 = 9'haf == r_count_9_io_out ? io_r_175_b : _GEN_3954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3956 = 9'hb0 == r_count_9_io_out ? io_r_176_b : _GEN_3955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3957 = 9'hb1 == r_count_9_io_out ? io_r_177_b : _GEN_3956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3958 = 9'hb2 == r_count_9_io_out ? io_r_178_b : _GEN_3957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3959 = 9'hb3 == r_count_9_io_out ? io_r_179_b : _GEN_3958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3960 = 9'hb4 == r_count_9_io_out ? io_r_180_b : _GEN_3959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3961 = 9'hb5 == r_count_9_io_out ? io_r_181_b : _GEN_3960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3962 = 9'hb6 == r_count_9_io_out ? io_r_182_b : _GEN_3961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3963 = 9'hb7 == r_count_9_io_out ? io_r_183_b : _GEN_3962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3964 = 9'hb8 == r_count_9_io_out ? io_r_184_b : _GEN_3963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3965 = 9'hb9 == r_count_9_io_out ? io_r_185_b : _GEN_3964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3966 = 9'hba == r_count_9_io_out ? io_r_186_b : _GEN_3965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3967 = 9'hbb == r_count_9_io_out ? io_r_187_b : _GEN_3966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3968 = 9'hbc == r_count_9_io_out ? io_r_188_b : _GEN_3967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3969 = 9'hbd == r_count_9_io_out ? io_r_189_b : _GEN_3968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3970 = 9'hbe == r_count_9_io_out ? io_r_190_b : _GEN_3969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3971 = 9'hbf == r_count_9_io_out ? io_r_191_b : _GEN_3970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3972 = 9'hc0 == r_count_9_io_out ? io_r_192_b : _GEN_3971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3973 = 9'hc1 == r_count_9_io_out ? io_r_193_b : _GEN_3972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3974 = 9'hc2 == r_count_9_io_out ? io_r_194_b : _GEN_3973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3975 = 9'hc3 == r_count_9_io_out ? io_r_195_b : _GEN_3974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3976 = 9'hc4 == r_count_9_io_out ? io_r_196_b : _GEN_3975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3977 = 9'hc5 == r_count_9_io_out ? io_r_197_b : _GEN_3976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3978 = 9'hc6 == r_count_9_io_out ? io_r_198_b : _GEN_3977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3979 = 9'hc7 == r_count_9_io_out ? io_r_199_b : _GEN_3978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3980 = 9'hc8 == r_count_9_io_out ? io_r_200_b : _GEN_3979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3981 = 9'hc9 == r_count_9_io_out ? io_r_201_b : _GEN_3980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3982 = 9'hca == r_count_9_io_out ? io_r_202_b : _GEN_3981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3983 = 9'hcb == r_count_9_io_out ? io_r_203_b : _GEN_3982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3984 = 9'hcc == r_count_9_io_out ? io_r_204_b : _GEN_3983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3985 = 9'hcd == r_count_9_io_out ? io_r_205_b : _GEN_3984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3986 = 9'hce == r_count_9_io_out ? io_r_206_b : _GEN_3985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3987 = 9'hcf == r_count_9_io_out ? io_r_207_b : _GEN_3986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3988 = 9'hd0 == r_count_9_io_out ? io_r_208_b : _GEN_3987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3989 = 9'hd1 == r_count_9_io_out ? io_r_209_b : _GEN_3988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3990 = 9'hd2 == r_count_9_io_out ? io_r_210_b : _GEN_3989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3991 = 9'hd3 == r_count_9_io_out ? io_r_211_b : _GEN_3990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3992 = 9'hd4 == r_count_9_io_out ? io_r_212_b : _GEN_3991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3993 = 9'hd5 == r_count_9_io_out ? io_r_213_b : _GEN_3992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3994 = 9'hd6 == r_count_9_io_out ? io_r_214_b : _GEN_3993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3995 = 9'hd7 == r_count_9_io_out ? io_r_215_b : _GEN_3994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3996 = 9'hd8 == r_count_9_io_out ? io_r_216_b : _GEN_3995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3997 = 9'hd9 == r_count_9_io_out ? io_r_217_b : _GEN_3996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3998 = 9'hda == r_count_9_io_out ? io_r_218_b : _GEN_3997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3999 = 9'hdb == r_count_9_io_out ? io_r_219_b : _GEN_3998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4000 = 9'hdc == r_count_9_io_out ? io_r_220_b : _GEN_3999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4001 = 9'hdd == r_count_9_io_out ? io_r_221_b : _GEN_4000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4002 = 9'hde == r_count_9_io_out ? io_r_222_b : _GEN_4001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4003 = 9'hdf == r_count_9_io_out ? io_r_223_b : _GEN_4002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4004 = 9'he0 == r_count_9_io_out ? io_r_224_b : _GEN_4003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4005 = 9'he1 == r_count_9_io_out ? io_r_225_b : _GEN_4004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4006 = 9'he2 == r_count_9_io_out ? io_r_226_b : _GEN_4005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4007 = 9'he3 == r_count_9_io_out ? io_r_227_b : _GEN_4006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4008 = 9'he4 == r_count_9_io_out ? io_r_228_b : _GEN_4007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4009 = 9'he5 == r_count_9_io_out ? io_r_229_b : _GEN_4008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4010 = 9'he6 == r_count_9_io_out ? io_r_230_b : _GEN_4009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4011 = 9'he7 == r_count_9_io_out ? io_r_231_b : _GEN_4010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4012 = 9'he8 == r_count_9_io_out ? io_r_232_b : _GEN_4011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4013 = 9'he9 == r_count_9_io_out ? io_r_233_b : _GEN_4012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4014 = 9'hea == r_count_9_io_out ? io_r_234_b : _GEN_4013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4015 = 9'heb == r_count_9_io_out ? io_r_235_b : _GEN_4014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4016 = 9'hec == r_count_9_io_out ? io_r_236_b : _GEN_4015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4017 = 9'hed == r_count_9_io_out ? io_r_237_b : _GEN_4016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4018 = 9'hee == r_count_9_io_out ? io_r_238_b : _GEN_4017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4019 = 9'hef == r_count_9_io_out ? io_r_239_b : _GEN_4018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4020 = 9'hf0 == r_count_9_io_out ? io_r_240_b : _GEN_4019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4021 = 9'hf1 == r_count_9_io_out ? io_r_241_b : _GEN_4020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4022 = 9'hf2 == r_count_9_io_out ? io_r_242_b : _GEN_4021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4023 = 9'hf3 == r_count_9_io_out ? io_r_243_b : _GEN_4022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4024 = 9'hf4 == r_count_9_io_out ? io_r_244_b : _GEN_4023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4025 = 9'hf5 == r_count_9_io_out ? io_r_245_b : _GEN_4024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4026 = 9'hf6 == r_count_9_io_out ? io_r_246_b : _GEN_4025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4027 = 9'hf7 == r_count_9_io_out ? io_r_247_b : _GEN_4026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4028 = 9'hf8 == r_count_9_io_out ? io_r_248_b : _GEN_4027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4029 = 9'hf9 == r_count_9_io_out ? io_r_249_b : _GEN_4028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4030 = 9'hfa == r_count_9_io_out ? io_r_250_b : _GEN_4029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4031 = 9'hfb == r_count_9_io_out ? io_r_251_b : _GEN_4030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4032 = 9'hfc == r_count_9_io_out ? io_r_252_b : _GEN_4031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4033 = 9'hfd == r_count_9_io_out ? io_r_253_b : _GEN_4032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4034 = 9'hfe == r_count_9_io_out ? io_r_254_b : _GEN_4033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4035 = 9'hff == r_count_9_io_out ? io_r_255_b : _GEN_4034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4036 = 9'h100 == r_count_9_io_out ? io_r_256_b : _GEN_4035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4037 = 9'h101 == r_count_9_io_out ? io_r_257_b : _GEN_4036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4038 = 9'h102 == r_count_9_io_out ? io_r_258_b : _GEN_4037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4039 = 9'h103 == r_count_9_io_out ? io_r_259_b : _GEN_4038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4040 = 9'h104 == r_count_9_io_out ? io_r_260_b : _GEN_4039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4041 = 9'h105 == r_count_9_io_out ? io_r_261_b : _GEN_4040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4042 = 9'h106 == r_count_9_io_out ? io_r_262_b : _GEN_4041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4043 = 9'h107 == r_count_9_io_out ? io_r_263_b : _GEN_4042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4044 = 9'h108 == r_count_9_io_out ? io_r_264_b : _GEN_4043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4045 = 9'h109 == r_count_9_io_out ? io_r_265_b : _GEN_4044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4046 = 9'h10a == r_count_9_io_out ? io_r_266_b : _GEN_4045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4047 = 9'h10b == r_count_9_io_out ? io_r_267_b : _GEN_4046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4048 = 9'h10c == r_count_9_io_out ? io_r_268_b : _GEN_4047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4049 = 9'h10d == r_count_9_io_out ? io_r_269_b : _GEN_4048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4050 = 9'h10e == r_count_9_io_out ? io_r_270_b : _GEN_4049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4051 = 9'h10f == r_count_9_io_out ? io_r_271_b : _GEN_4050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4052 = 9'h110 == r_count_9_io_out ? io_r_272_b : _GEN_4051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4053 = 9'h111 == r_count_9_io_out ? io_r_273_b : _GEN_4052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4054 = 9'h112 == r_count_9_io_out ? io_r_274_b : _GEN_4053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4055 = 9'h113 == r_count_9_io_out ? io_r_275_b : _GEN_4054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4056 = 9'h114 == r_count_9_io_out ? io_r_276_b : _GEN_4055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4057 = 9'h115 == r_count_9_io_out ? io_r_277_b : _GEN_4056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4058 = 9'h116 == r_count_9_io_out ? io_r_278_b : _GEN_4057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4059 = 9'h117 == r_count_9_io_out ? io_r_279_b : _GEN_4058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4060 = 9'h118 == r_count_9_io_out ? io_r_280_b : _GEN_4059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4061 = 9'h119 == r_count_9_io_out ? io_r_281_b : _GEN_4060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4062 = 9'h11a == r_count_9_io_out ? io_r_282_b : _GEN_4061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4063 = 9'h11b == r_count_9_io_out ? io_r_283_b : _GEN_4062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4064 = 9'h11c == r_count_9_io_out ? io_r_284_b : _GEN_4063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4065 = 9'h11d == r_count_9_io_out ? io_r_285_b : _GEN_4064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4066 = 9'h11e == r_count_9_io_out ? io_r_286_b : _GEN_4065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4067 = 9'h11f == r_count_9_io_out ? io_r_287_b : _GEN_4066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4068 = 9'h120 == r_count_9_io_out ? io_r_288_b : _GEN_4067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4069 = 9'h121 == r_count_9_io_out ? io_r_289_b : _GEN_4068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4070 = 9'h122 == r_count_9_io_out ? io_r_290_b : _GEN_4069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4071 = 9'h123 == r_count_9_io_out ? io_r_291_b : _GEN_4070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4072 = 9'h124 == r_count_9_io_out ? io_r_292_b : _GEN_4071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4073 = 9'h125 == r_count_9_io_out ? io_r_293_b : _GEN_4072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4074 = 9'h126 == r_count_9_io_out ? io_r_294_b : _GEN_4073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4075 = 9'h127 == r_count_9_io_out ? io_r_295_b : _GEN_4074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4076 = 9'h128 == r_count_9_io_out ? io_r_296_b : _GEN_4075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4077 = 9'h129 == r_count_9_io_out ? io_r_297_b : _GEN_4076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4078 = 9'h12a == r_count_9_io_out ? io_r_298_b : _GEN_4077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4079 = 9'h12b == r_count_9_io_out ? io_r_299_b : _GEN_4078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4080 = 9'h12c == r_count_9_io_out ? io_r_300_b : _GEN_4079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4081 = 9'h12d == r_count_9_io_out ? io_r_301_b : _GEN_4080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4082 = 9'h12e == r_count_9_io_out ? io_r_302_b : _GEN_4081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4083 = 9'h12f == r_count_9_io_out ? io_r_303_b : _GEN_4082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4084 = 9'h130 == r_count_9_io_out ? io_r_304_b : _GEN_4083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4085 = 9'h131 == r_count_9_io_out ? io_r_305_b : _GEN_4084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4086 = 9'h132 == r_count_9_io_out ? io_r_306_b : _GEN_4085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4087 = 9'h133 == r_count_9_io_out ? io_r_307_b : _GEN_4086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4088 = 9'h134 == r_count_9_io_out ? io_r_308_b : _GEN_4087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4089 = 9'h135 == r_count_9_io_out ? io_r_309_b : _GEN_4088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4090 = 9'h136 == r_count_9_io_out ? io_r_310_b : _GEN_4089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4091 = 9'h137 == r_count_9_io_out ? io_r_311_b : _GEN_4090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4092 = 9'h138 == r_count_9_io_out ? io_r_312_b : _GEN_4091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4093 = 9'h139 == r_count_9_io_out ? io_r_313_b : _GEN_4092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4094 = 9'h13a == r_count_9_io_out ? io_r_314_b : _GEN_4093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4095 = 9'h13b == r_count_9_io_out ? io_r_315_b : _GEN_4094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4096 = 9'h13c == r_count_9_io_out ? io_r_316_b : _GEN_4095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4097 = 9'h13d == r_count_9_io_out ? io_r_317_b : _GEN_4096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4098 = 9'h13e == r_count_9_io_out ? io_r_318_b : _GEN_4097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4099 = 9'h13f == r_count_9_io_out ? io_r_319_b : _GEN_4098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4100 = 9'h140 == r_count_9_io_out ? io_r_320_b : _GEN_4099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4101 = 9'h141 == r_count_9_io_out ? io_r_321_b : _GEN_4100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4102 = 9'h142 == r_count_9_io_out ? io_r_322_b : _GEN_4101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4103 = 9'h143 == r_count_9_io_out ? io_r_323_b : _GEN_4102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4104 = 9'h144 == r_count_9_io_out ? io_r_324_b : _GEN_4103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4105 = 9'h145 == r_count_9_io_out ? io_r_325_b : _GEN_4104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4106 = 9'h146 == r_count_9_io_out ? io_r_326_b : _GEN_4105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4107 = 9'h147 == r_count_9_io_out ? io_r_327_b : _GEN_4106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4108 = 9'h148 == r_count_9_io_out ? io_r_328_b : _GEN_4107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4109 = 9'h149 == r_count_9_io_out ? io_r_329_b : _GEN_4108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4110 = 9'h14a == r_count_9_io_out ? io_r_330_b : _GEN_4109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4111 = 9'h14b == r_count_9_io_out ? io_r_331_b : _GEN_4110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4112 = 9'h14c == r_count_9_io_out ? io_r_332_b : _GEN_4111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4113 = 9'h14d == r_count_9_io_out ? io_r_333_b : _GEN_4112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4114 = 9'h14e == r_count_9_io_out ? io_r_334_b : _GEN_4113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4115 = 9'h14f == r_count_9_io_out ? io_r_335_b : _GEN_4114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4116 = 9'h150 == r_count_9_io_out ? io_r_336_b : _GEN_4115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4117 = 9'h151 == r_count_9_io_out ? io_r_337_b : _GEN_4116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4118 = 9'h152 == r_count_9_io_out ? io_r_338_b : _GEN_4117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4119 = 9'h153 == r_count_9_io_out ? io_r_339_b : _GEN_4118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4120 = 9'h154 == r_count_9_io_out ? io_r_340_b : _GEN_4119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4121 = 9'h155 == r_count_9_io_out ? io_r_341_b : _GEN_4120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4122 = 9'h156 == r_count_9_io_out ? io_r_342_b : _GEN_4121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4123 = 9'h157 == r_count_9_io_out ? io_r_343_b : _GEN_4122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4124 = 9'h158 == r_count_9_io_out ? io_r_344_b : _GEN_4123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4125 = 9'h159 == r_count_9_io_out ? io_r_345_b : _GEN_4124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4126 = 9'h15a == r_count_9_io_out ? io_r_346_b : _GEN_4125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4127 = 9'h15b == r_count_9_io_out ? io_r_347_b : _GEN_4126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4128 = 9'h15c == r_count_9_io_out ? io_r_348_b : _GEN_4127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4129 = 9'h15d == r_count_9_io_out ? io_r_349_b : _GEN_4128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4130 = 9'h15e == r_count_9_io_out ? io_r_350_b : _GEN_4129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4131 = 9'h15f == r_count_9_io_out ? io_r_351_b : _GEN_4130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4132 = 9'h160 == r_count_9_io_out ? io_r_352_b : _GEN_4131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4133 = 9'h161 == r_count_9_io_out ? io_r_353_b : _GEN_4132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4134 = 9'h162 == r_count_9_io_out ? io_r_354_b : _GEN_4133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4135 = 9'h163 == r_count_9_io_out ? io_r_355_b : _GEN_4134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4136 = 9'h164 == r_count_9_io_out ? io_r_356_b : _GEN_4135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4137 = 9'h165 == r_count_9_io_out ? io_r_357_b : _GEN_4136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4138 = 9'h166 == r_count_9_io_out ? io_r_358_b : _GEN_4137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4139 = 9'h167 == r_count_9_io_out ? io_r_359_b : _GEN_4138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4140 = 9'h168 == r_count_9_io_out ? io_r_360_b : _GEN_4139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4141 = 9'h169 == r_count_9_io_out ? io_r_361_b : _GEN_4140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4142 = 9'h16a == r_count_9_io_out ? io_r_362_b : _GEN_4141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4143 = 9'h16b == r_count_9_io_out ? io_r_363_b : _GEN_4142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4144 = 9'h16c == r_count_9_io_out ? io_r_364_b : _GEN_4143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4145 = 9'h16d == r_count_9_io_out ? io_r_365_b : _GEN_4144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4146 = 9'h16e == r_count_9_io_out ? io_r_366_b : _GEN_4145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4147 = 9'h16f == r_count_9_io_out ? io_r_367_b : _GEN_4146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4148 = 9'h170 == r_count_9_io_out ? io_r_368_b : _GEN_4147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4149 = 9'h171 == r_count_9_io_out ? io_r_369_b : _GEN_4148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4150 = 9'h172 == r_count_9_io_out ? io_r_370_b : _GEN_4149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4151 = 9'h173 == r_count_9_io_out ? io_r_371_b : _GEN_4150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4152 = 9'h174 == r_count_9_io_out ? io_r_372_b : _GEN_4151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4153 = 9'h175 == r_count_9_io_out ? io_r_373_b : _GEN_4152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4154 = 9'h176 == r_count_9_io_out ? io_r_374_b : _GEN_4153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4155 = 9'h177 == r_count_9_io_out ? io_r_375_b : _GEN_4154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4156 = 9'h178 == r_count_9_io_out ? io_r_376_b : _GEN_4155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4157 = 9'h179 == r_count_9_io_out ? io_r_377_b : _GEN_4156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4158 = 9'h17a == r_count_9_io_out ? io_r_378_b : _GEN_4157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4159 = 9'h17b == r_count_9_io_out ? io_r_379_b : _GEN_4158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4160 = 9'h17c == r_count_9_io_out ? io_r_380_b : _GEN_4159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4161 = 9'h17d == r_count_9_io_out ? io_r_381_b : _GEN_4160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4162 = 9'h17e == r_count_9_io_out ? io_r_382_b : _GEN_4161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4163 = 9'h17f == r_count_9_io_out ? io_r_383_b : _GEN_4162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4164 = 9'h180 == r_count_9_io_out ? io_r_384_b : _GEN_4163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4165 = 9'h181 == r_count_9_io_out ? io_r_385_b : _GEN_4164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4166 = 9'h182 == r_count_9_io_out ? io_r_386_b : _GEN_4165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4167 = 9'h183 == r_count_9_io_out ? io_r_387_b : _GEN_4166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4168 = 9'h184 == r_count_9_io_out ? io_r_388_b : _GEN_4167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4169 = 9'h185 == r_count_9_io_out ? io_r_389_b : _GEN_4168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4170 = 9'h186 == r_count_9_io_out ? io_r_390_b : _GEN_4169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4171 = 9'h187 == r_count_9_io_out ? io_r_391_b : _GEN_4170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4172 = 9'h188 == r_count_9_io_out ? io_r_392_b : _GEN_4171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4173 = 9'h189 == r_count_9_io_out ? io_r_393_b : _GEN_4172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4174 = 9'h18a == r_count_9_io_out ? io_r_394_b : _GEN_4173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4175 = 9'h18b == r_count_9_io_out ? io_r_395_b : _GEN_4174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4176 = 9'h18c == r_count_9_io_out ? io_r_396_b : _GEN_4175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4177 = 9'h18d == r_count_9_io_out ? io_r_397_b : _GEN_4176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4178 = 9'h18e == r_count_9_io_out ? io_r_398_b : _GEN_4177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4181 = 9'h1 == r_count_10_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4182 = 9'h2 == r_count_10_io_out ? io_r_2_b : _GEN_4181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4183 = 9'h3 == r_count_10_io_out ? io_r_3_b : _GEN_4182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4184 = 9'h4 == r_count_10_io_out ? io_r_4_b : _GEN_4183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4185 = 9'h5 == r_count_10_io_out ? io_r_5_b : _GEN_4184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4186 = 9'h6 == r_count_10_io_out ? io_r_6_b : _GEN_4185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4187 = 9'h7 == r_count_10_io_out ? io_r_7_b : _GEN_4186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4188 = 9'h8 == r_count_10_io_out ? io_r_8_b : _GEN_4187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4189 = 9'h9 == r_count_10_io_out ? io_r_9_b : _GEN_4188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4190 = 9'ha == r_count_10_io_out ? io_r_10_b : _GEN_4189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4191 = 9'hb == r_count_10_io_out ? io_r_11_b : _GEN_4190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4192 = 9'hc == r_count_10_io_out ? io_r_12_b : _GEN_4191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4193 = 9'hd == r_count_10_io_out ? io_r_13_b : _GEN_4192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4194 = 9'he == r_count_10_io_out ? io_r_14_b : _GEN_4193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4195 = 9'hf == r_count_10_io_out ? io_r_15_b : _GEN_4194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4196 = 9'h10 == r_count_10_io_out ? io_r_16_b : _GEN_4195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4197 = 9'h11 == r_count_10_io_out ? io_r_17_b : _GEN_4196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4198 = 9'h12 == r_count_10_io_out ? io_r_18_b : _GEN_4197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4199 = 9'h13 == r_count_10_io_out ? io_r_19_b : _GEN_4198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4200 = 9'h14 == r_count_10_io_out ? io_r_20_b : _GEN_4199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4201 = 9'h15 == r_count_10_io_out ? io_r_21_b : _GEN_4200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4202 = 9'h16 == r_count_10_io_out ? io_r_22_b : _GEN_4201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4203 = 9'h17 == r_count_10_io_out ? io_r_23_b : _GEN_4202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4204 = 9'h18 == r_count_10_io_out ? io_r_24_b : _GEN_4203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4205 = 9'h19 == r_count_10_io_out ? io_r_25_b : _GEN_4204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4206 = 9'h1a == r_count_10_io_out ? io_r_26_b : _GEN_4205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4207 = 9'h1b == r_count_10_io_out ? io_r_27_b : _GEN_4206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4208 = 9'h1c == r_count_10_io_out ? io_r_28_b : _GEN_4207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4209 = 9'h1d == r_count_10_io_out ? io_r_29_b : _GEN_4208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4210 = 9'h1e == r_count_10_io_out ? io_r_30_b : _GEN_4209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4211 = 9'h1f == r_count_10_io_out ? io_r_31_b : _GEN_4210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4212 = 9'h20 == r_count_10_io_out ? io_r_32_b : _GEN_4211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4213 = 9'h21 == r_count_10_io_out ? io_r_33_b : _GEN_4212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4214 = 9'h22 == r_count_10_io_out ? io_r_34_b : _GEN_4213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4215 = 9'h23 == r_count_10_io_out ? io_r_35_b : _GEN_4214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4216 = 9'h24 == r_count_10_io_out ? io_r_36_b : _GEN_4215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4217 = 9'h25 == r_count_10_io_out ? io_r_37_b : _GEN_4216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4218 = 9'h26 == r_count_10_io_out ? io_r_38_b : _GEN_4217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4219 = 9'h27 == r_count_10_io_out ? io_r_39_b : _GEN_4218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4220 = 9'h28 == r_count_10_io_out ? io_r_40_b : _GEN_4219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4221 = 9'h29 == r_count_10_io_out ? io_r_41_b : _GEN_4220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4222 = 9'h2a == r_count_10_io_out ? io_r_42_b : _GEN_4221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4223 = 9'h2b == r_count_10_io_out ? io_r_43_b : _GEN_4222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4224 = 9'h2c == r_count_10_io_out ? io_r_44_b : _GEN_4223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4225 = 9'h2d == r_count_10_io_out ? io_r_45_b : _GEN_4224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4226 = 9'h2e == r_count_10_io_out ? io_r_46_b : _GEN_4225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4227 = 9'h2f == r_count_10_io_out ? io_r_47_b : _GEN_4226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4228 = 9'h30 == r_count_10_io_out ? io_r_48_b : _GEN_4227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4229 = 9'h31 == r_count_10_io_out ? io_r_49_b : _GEN_4228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4230 = 9'h32 == r_count_10_io_out ? io_r_50_b : _GEN_4229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4231 = 9'h33 == r_count_10_io_out ? io_r_51_b : _GEN_4230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4232 = 9'h34 == r_count_10_io_out ? io_r_52_b : _GEN_4231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4233 = 9'h35 == r_count_10_io_out ? io_r_53_b : _GEN_4232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4234 = 9'h36 == r_count_10_io_out ? io_r_54_b : _GEN_4233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4235 = 9'h37 == r_count_10_io_out ? io_r_55_b : _GEN_4234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4236 = 9'h38 == r_count_10_io_out ? io_r_56_b : _GEN_4235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4237 = 9'h39 == r_count_10_io_out ? io_r_57_b : _GEN_4236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4238 = 9'h3a == r_count_10_io_out ? io_r_58_b : _GEN_4237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4239 = 9'h3b == r_count_10_io_out ? io_r_59_b : _GEN_4238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4240 = 9'h3c == r_count_10_io_out ? io_r_60_b : _GEN_4239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4241 = 9'h3d == r_count_10_io_out ? io_r_61_b : _GEN_4240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4242 = 9'h3e == r_count_10_io_out ? io_r_62_b : _GEN_4241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4243 = 9'h3f == r_count_10_io_out ? io_r_63_b : _GEN_4242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4244 = 9'h40 == r_count_10_io_out ? io_r_64_b : _GEN_4243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4245 = 9'h41 == r_count_10_io_out ? io_r_65_b : _GEN_4244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4246 = 9'h42 == r_count_10_io_out ? io_r_66_b : _GEN_4245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4247 = 9'h43 == r_count_10_io_out ? io_r_67_b : _GEN_4246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4248 = 9'h44 == r_count_10_io_out ? io_r_68_b : _GEN_4247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4249 = 9'h45 == r_count_10_io_out ? io_r_69_b : _GEN_4248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4250 = 9'h46 == r_count_10_io_out ? io_r_70_b : _GEN_4249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4251 = 9'h47 == r_count_10_io_out ? io_r_71_b : _GEN_4250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4252 = 9'h48 == r_count_10_io_out ? io_r_72_b : _GEN_4251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4253 = 9'h49 == r_count_10_io_out ? io_r_73_b : _GEN_4252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4254 = 9'h4a == r_count_10_io_out ? io_r_74_b : _GEN_4253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4255 = 9'h4b == r_count_10_io_out ? io_r_75_b : _GEN_4254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4256 = 9'h4c == r_count_10_io_out ? io_r_76_b : _GEN_4255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4257 = 9'h4d == r_count_10_io_out ? io_r_77_b : _GEN_4256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4258 = 9'h4e == r_count_10_io_out ? io_r_78_b : _GEN_4257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4259 = 9'h4f == r_count_10_io_out ? io_r_79_b : _GEN_4258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4260 = 9'h50 == r_count_10_io_out ? io_r_80_b : _GEN_4259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4261 = 9'h51 == r_count_10_io_out ? io_r_81_b : _GEN_4260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4262 = 9'h52 == r_count_10_io_out ? io_r_82_b : _GEN_4261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4263 = 9'h53 == r_count_10_io_out ? io_r_83_b : _GEN_4262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4264 = 9'h54 == r_count_10_io_out ? io_r_84_b : _GEN_4263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4265 = 9'h55 == r_count_10_io_out ? io_r_85_b : _GEN_4264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4266 = 9'h56 == r_count_10_io_out ? io_r_86_b : _GEN_4265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4267 = 9'h57 == r_count_10_io_out ? io_r_87_b : _GEN_4266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4268 = 9'h58 == r_count_10_io_out ? io_r_88_b : _GEN_4267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4269 = 9'h59 == r_count_10_io_out ? io_r_89_b : _GEN_4268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4270 = 9'h5a == r_count_10_io_out ? io_r_90_b : _GEN_4269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4271 = 9'h5b == r_count_10_io_out ? io_r_91_b : _GEN_4270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4272 = 9'h5c == r_count_10_io_out ? io_r_92_b : _GEN_4271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4273 = 9'h5d == r_count_10_io_out ? io_r_93_b : _GEN_4272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4274 = 9'h5e == r_count_10_io_out ? io_r_94_b : _GEN_4273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4275 = 9'h5f == r_count_10_io_out ? io_r_95_b : _GEN_4274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4276 = 9'h60 == r_count_10_io_out ? io_r_96_b : _GEN_4275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4277 = 9'h61 == r_count_10_io_out ? io_r_97_b : _GEN_4276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4278 = 9'h62 == r_count_10_io_out ? io_r_98_b : _GEN_4277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4279 = 9'h63 == r_count_10_io_out ? io_r_99_b : _GEN_4278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4280 = 9'h64 == r_count_10_io_out ? io_r_100_b : _GEN_4279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4281 = 9'h65 == r_count_10_io_out ? io_r_101_b : _GEN_4280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4282 = 9'h66 == r_count_10_io_out ? io_r_102_b : _GEN_4281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4283 = 9'h67 == r_count_10_io_out ? io_r_103_b : _GEN_4282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4284 = 9'h68 == r_count_10_io_out ? io_r_104_b : _GEN_4283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4285 = 9'h69 == r_count_10_io_out ? io_r_105_b : _GEN_4284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4286 = 9'h6a == r_count_10_io_out ? io_r_106_b : _GEN_4285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4287 = 9'h6b == r_count_10_io_out ? io_r_107_b : _GEN_4286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4288 = 9'h6c == r_count_10_io_out ? io_r_108_b : _GEN_4287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4289 = 9'h6d == r_count_10_io_out ? io_r_109_b : _GEN_4288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4290 = 9'h6e == r_count_10_io_out ? io_r_110_b : _GEN_4289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4291 = 9'h6f == r_count_10_io_out ? io_r_111_b : _GEN_4290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4292 = 9'h70 == r_count_10_io_out ? io_r_112_b : _GEN_4291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4293 = 9'h71 == r_count_10_io_out ? io_r_113_b : _GEN_4292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4294 = 9'h72 == r_count_10_io_out ? io_r_114_b : _GEN_4293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4295 = 9'h73 == r_count_10_io_out ? io_r_115_b : _GEN_4294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4296 = 9'h74 == r_count_10_io_out ? io_r_116_b : _GEN_4295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4297 = 9'h75 == r_count_10_io_out ? io_r_117_b : _GEN_4296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4298 = 9'h76 == r_count_10_io_out ? io_r_118_b : _GEN_4297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4299 = 9'h77 == r_count_10_io_out ? io_r_119_b : _GEN_4298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4300 = 9'h78 == r_count_10_io_out ? io_r_120_b : _GEN_4299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4301 = 9'h79 == r_count_10_io_out ? io_r_121_b : _GEN_4300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4302 = 9'h7a == r_count_10_io_out ? io_r_122_b : _GEN_4301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4303 = 9'h7b == r_count_10_io_out ? io_r_123_b : _GEN_4302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4304 = 9'h7c == r_count_10_io_out ? io_r_124_b : _GEN_4303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4305 = 9'h7d == r_count_10_io_out ? io_r_125_b : _GEN_4304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4306 = 9'h7e == r_count_10_io_out ? io_r_126_b : _GEN_4305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4307 = 9'h7f == r_count_10_io_out ? io_r_127_b : _GEN_4306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4308 = 9'h80 == r_count_10_io_out ? io_r_128_b : _GEN_4307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4309 = 9'h81 == r_count_10_io_out ? io_r_129_b : _GEN_4308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4310 = 9'h82 == r_count_10_io_out ? io_r_130_b : _GEN_4309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4311 = 9'h83 == r_count_10_io_out ? io_r_131_b : _GEN_4310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4312 = 9'h84 == r_count_10_io_out ? io_r_132_b : _GEN_4311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4313 = 9'h85 == r_count_10_io_out ? io_r_133_b : _GEN_4312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4314 = 9'h86 == r_count_10_io_out ? io_r_134_b : _GEN_4313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4315 = 9'h87 == r_count_10_io_out ? io_r_135_b : _GEN_4314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4316 = 9'h88 == r_count_10_io_out ? io_r_136_b : _GEN_4315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4317 = 9'h89 == r_count_10_io_out ? io_r_137_b : _GEN_4316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4318 = 9'h8a == r_count_10_io_out ? io_r_138_b : _GEN_4317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4319 = 9'h8b == r_count_10_io_out ? io_r_139_b : _GEN_4318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4320 = 9'h8c == r_count_10_io_out ? io_r_140_b : _GEN_4319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4321 = 9'h8d == r_count_10_io_out ? io_r_141_b : _GEN_4320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4322 = 9'h8e == r_count_10_io_out ? io_r_142_b : _GEN_4321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4323 = 9'h8f == r_count_10_io_out ? io_r_143_b : _GEN_4322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4324 = 9'h90 == r_count_10_io_out ? io_r_144_b : _GEN_4323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4325 = 9'h91 == r_count_10_io_out ? io_r_145_b : _GEN_4324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4326 = 9'h92 == r_count_10_io_out ? io_r_146_b : _GEN_4325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4327 = 9'h93 == r_count_10_io_out ? io_r_147_b : _GEN_4326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4328 = 9'h94 == r_count_10_io_out ? io_r_148_b : _GEN_4327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4329 = 9'h95 == r_count_10_io_out ? io_r_149_b : _GEN_4328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4330 = 9'h96 == r_count_10_io_out ? io_r_150_b : _GEN_4329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4331 = 9'h97 == r_count_10_io_out ? io_r_151_b : _GEN_4330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4332 = 9'h98 == r_count_10_io_out ? io_r_152_b : _GEN_4331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4333 = 9'h99 == r_count_10_io_out ? io_r_153_b : _GEN_4332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4334 = 9'h9a == r_count_10_io_out ? io_r_154_b : _GEN_4333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4335 = 9'h9b == r_count_10_io_out ? io_r_155_b : _GEN_4334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4336 = 9'h9c == r_count_10_io_out ? io_r_156_b : _GEN_4335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4337 = 9'h9d == r_count_10_io_out ? io_r_157_b : _GEN_4336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4338 = 9'h9e == r_count_10_io_out ? io_r_158_b : _GEN_4337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4339 = 9'h9f == r_count_10_io_out ? io_r_159_b : _GEN_4338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4340 = 9'ha0 == r_count_10_io_out ? io_r_160_b : _GEN_4339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4341 = 9'ha1 == r_count_10_io_out ? io_r_161_b : _GEN_4340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4342 = 9'ha2 == r_count_10_io_out ? io_r_162_b : _GEN_4341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4343 = 9'ha3 == r_count_10_io_out ? io_r_163_b : _GEN_4342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4344 = 9'ha4 == r_count_10_io_out ? io_r_164_b : _GEN_4343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4345 = 9'ha5 == r_count_10_io_out ? io_r_165_b : _GEN_4344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4346 = 9'ha6 == r_count_10_io_out ? io_r_166_b : _GEN_4345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4347 = 9'ha7 == r_count_10_io_out ? io_r_167_b : _GEN_4346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4348 = 9'ha8 == r_count_10_io_out ? io_r_168_b : _GEN_4347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4349 = 9'ha9 == r_count_10_io_out ? io_r_169_b : _GEN_4348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4350 = 9'haa == r_count_10_io_out ? io_r_170_b : _GEN_4349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4351 = 9'hab == r_count_10_io_out ? io_r_171_b : _GEN_4350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4352 = 9'hac == r_count_10_io_out ? io_r_172_b : _GEN_4351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4353 = 9'had == r_count_10_io_out ? io_r_173_b : _GEN_4352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4354 = 9'hae == r_count_10_io_out ? io_r_174_b : _GEN_4353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4355 = 9'haf == r_count_10_io_out ? io_r_175_b : _GEN_4354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4356 = 9'hb0 == r_count_10_io_out ? io_r_176_b : _GEN_4355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4357 = 9'hb1 == r_count_10_io_out ? io_r_177_b : _GEN_4356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4358 = 9'hb2 == r_count_10_io_out ? io_r_178_b : _GEN_4357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4359 = 9'hb3 == r_count_10_io_out ? io_r_179_b : _GEN_4358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4360 = 9'hb4 == r_count_10_io_out ? io_r_180_b : _GEN_4359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4361 = 9'hb5 == r_count_10_io_out ? io_r_181_b : _GEN_4360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4362 = 9'hb6 == r_count_10_io_out ? io_r_182_b : _GEN_4361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4363 = 9'hb7 == r_count_10_io_out ? io_r_183_b : _GEN_4362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4364 = 9'hb8 == r_count_10_io_out ? io_r_184_b : _GEN_4363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4365 = 9'hb9 == r_count_10_io_out ? io_r_185_b : _GEN_4364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4366 = 9'hba == r_count_10_io_out ? io_r_186_b : _GEN_4365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4367 = 9'hbb == r_count_10_io_out ? io_r_187_b : _GEN_4366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4368 = 9'hbc == r_count_10_io_out ? io_r_188_b : _GEN_4367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4369 = 9'hbd == r_count_10_io_out ? io_r_189_b : _GEN_4368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4370 = 9'hbe == r_count_10_io_out ? io_r_190_b : _GEN_4369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4371 = 9'hbf == r_count_10_io_out ? io_r_191_b : _GEN_4370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4372 = 9'hc0 == r_count_10_io_out ? io_r_192_b : _GEN_4371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4373 = 9'hc1 == r_count_10_io_out ? io_r_193_b : _GEN_4372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4374 = 9'hc2 == r_count_10_io_out ? io_r_194_b : _GEN_4373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4375 = 9'hc3 == r_count_10_io_out ? io_r_195_b : _GEN_4374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4376 = 9'hc4 == r_count_10_io_out ? io_r_196_b : _GEN_4375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4377 = 9'hc5 == r_count_10_io_out ? io_r_197_b : _GEN_4376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4378 = 9'hc6 == r_count_10_io_out ? io_r_198_b : _GEN_4377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4379 = 9'hc7 == r_count_10_io_out ? io_r_199_b : _GEN_4378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4380 = 9'hc8 == r_count_10_io_out ? io_r_200_b : _GEN_4379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4381 = 9'hc9 == r_count_10_io_out ? io_r_201_b : _GEN_4380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4382 = 9'hca == r_count_10_io_out ? io_r_202_b : _GEN_4381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4383 = 9'hcb == r_count_10_io_out ? io_r_203_b : _GEN_4382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4384 = 9'hcc == r_count_10_io_out ? io_r_204_b : _GEN_4383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4385 = 9'hcd == r_count_10_io_out ? io_r_205_b : _GEN_4384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4386 = 9'hce == r_count_10_io_out ? io_r_206_b : _GEN_4385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4387 = 9'hcf == r_count_10_io_out ? io_r_207_b : _GEN_4386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4388 = 9'hd0 == r_count_10_io_out ? io_r_208_b : _GEN_4387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4389 = 9'hd1 == r_count_10_io_out ? io_r_209_b : _GEN_4388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4390 = 9'hd2 == r_count_10_io_out ? io_r_210_b : _GEN_4389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4391 = 9'hd3 == r_count_10_io_out ? io_r_211_b : _GEN_4390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4392 = 9'hd4 == r_count_10_io_out ? io_r_212_b : _GEN_4391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4393 = 9'hd5 == r_count_10_io_out ? io_r_213_b : _GEN_4392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4394 = 9'hd6 == r_count_10_io_out ? io_r_214_b : _GEN_4393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4395 = 9'hd7 == r_count_10_io_out ? io_r_215_b : _GEN_4394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4396 = 9'hd8 == r_count_10_io_out ? io_r_216_b : _GEN_4395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4397 = 9'hd9 == r_count_10_io_out ? io_r_217_b : _GEN_4396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4398 = 9'hda == r_count_10_io_out ? io_r_218_b : _GEN_4397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4399 = 9'hdb == r_count_10_io_out ? io_r_219_b : _GEN_4398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4400 = 9'hdc == r_count_10_io_out ? io_r_220_b : _GEN_4399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4401 = 9'hdd == r_count_10_io_out ? io_r_221_b : _GEN_4400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4402 = 9'hde == r_count_10_io_out ? io_r_222_b : _GEN_4401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4403 = 9'hdf == r_count_10_io_out ? io_r_223_b : _GEN_4402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4404 = 9'he0 == r_count_10_io_out ? io_r_224_b : _GEN_4403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4405 = 9'he1 == r_count_10_io_out ? io_r_225_b : _GEN_4404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4406 = 9'he2 == r_count_10_io_out ? io_r_226_b : _GEN_4405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4407 = 9'he3 == r_count_10_io_out ? io_r_227_b : _GEN_4406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4408 = 9'he4 == r_count_10_io_out ? io_r_228_b : _GEN_4407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4409 = 9'he5 == r_count_10_io_out ? io_r_229_b : _GEN_4408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4410 = 9'he6 == r_count_10_io_out ? io_r_230_b : _GEN_4409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4411 = 9'he7 == r_count_10_io_out ? io_r_231_b : _GEN_4410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4412 = 9'he8 == r_count_10_io_out ? io_r_232_b : _GEN_4411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4413 = 9'he9 == r_count_10_io_out ? io_r_233_b : _GEN_4412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4414 = 9'hea == r_count_10_io_out ? io_r_234_b : _GEN_4413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4415 = 9'heb == r_count_10_io_out ? io_r_235_b : _GEN_4414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4416 = 9'hec == r_count_10_io_out ? io_r_236_b : _GEN_4415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4417 = 9'hed == r_count_10_io_out ? io_r_237_b : _GEN_4416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4418 = 9'hee == r_count_10_io_out ? io_r_238_b : _GEN_4417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4419 = 9'hef == r_count_10_io_out ? io_r_239_b : _GEN_4418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4420 = 9'hf0 == r_count_10_io_out ? io_r_240_b : _GEN_4419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4421 = 9'hf1 == r_count_10_io_out ? io_r_241_b : _GEN_4420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4422 = 9'hf2 == r_count_10_io_out ? io_r_242_b : _GEN_4421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4423 = 9'hf3 == r_count_10_io_out ? io_r_243_b : _GEN_4422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4424 = 9'hf4 == r_count_10_io_out ? io_r_244_b : _GEN_4423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4425 = 9'hf5 == r_count_10_io_out ? io_r_245_b : _GEN_4424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4426 = 9'hf6 == r_count_10_io_out ? io_r_246_b : _GEN_4425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4427 = 9'hf7 == r_count_10_io_out ? io_r_247_b : _GEN_4426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4428 = 9'hf8 == r_count_10_io_out ? io_r_248_b : _GEN_4427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4429 = 9'hf9 == r_count_10_io_out ? io_r_249_b : _GEN_4428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4430 = 9'hfa == r_count_10_io_out ? io_r_250_b : _GEN_4429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4431 = 9'hfb == r_count_10_io_out ? io_r_251_b : _GEN_4430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4432 = 9'hfc == r_count_10_io_out ? io_r_252_b : _GEN_4431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4433 = 9'hfd == r_count_10_io_out ? io_r_253_b : _GEN_4432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4434 = 9'hfe == r_count_10_io_out ? io_r_254_b : _GEN_4433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4435 = 9'hff == r_count_10_io_out ? io_r_255_b : _GEN_4434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4436 = 9'h100 == r_count_10_io_out ? io_r_256_b : _GEN_4435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4437 = 9'h101 == r_count_10_io_out ? io_r_257_b : _GEN_4436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4438 = 9'h102 == r_count_10_io_out ? io_r_258_b : _GEN_4437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4439 = 9'h103 == r_count_10_io_out ? io_r_259_b : _GEN_4438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4440 = 9'h104 == r_count_10_io_out ? io_r_260_b : _GEN_4439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4441 = 9'h105 == r_count_10_io_out ? io_r_261_b : _GEN_4440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4442 = 9'h106 == r_count_10_io_out ? io_r_262_b : _GEN_4441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4443 = 9'h107 == r_count_10_io_out ? io_r_263_b : _GEN_4442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4444 = 9'h108 == r_count_10_io_out ? io_r_264_b : _GEN_4443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4445 = 9'h109 == r_count_10_io_out ? io_r_265_b : _GEN_4444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4446 = 9'h10a == r_count_10_io_out ? io_r_266_b : _GEN_4445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4447 = 9'h10b == r_count_10_io_out ? io_r_267_b : _GEN_4446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4448 = 9'h10c == r_count_10_io_out ? io_r_268_b : _GEN_4447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4449 = 9'h10d == r_count_10_io_out ? io_r_269_b : _GEN_4448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4450 = 9'h10e == r_count_10_io_out ? io_r_270_b : _GEN_4449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4451 = 9'h10f == r_count_10_io_out ? io_r_271_b : _GEN_4450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4452 = 9'h110 == r_count_10_io_out ? io_r_272_b : _GEN_4451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4453 = 9'h111 == r_count_10_io_out ? io_r_273_b : _GEN_4452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4454 = 9'h112 == r_count_10_io_out ? io_r_274_b : _GEN_4453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4455 = 9'h113 == r_count_10_io_out ? io_r_275_b : _GEN_4454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4456 = 9'h114 == r_count_10_io_out ? io_r_276_b : _GEN_4455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4457 = 9'h115 == r_count_10_io_out ? io_r_277_b : _GEN_4456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4458 = 9'h116 == r_count_10_io_out ? io_r_278_b : _GEN_4457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4459 = 9'h117 == r_count_10_io_out ? io_r_279_b : _GEN_4458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4460 = 9'h118 == r_count_10_io_out ? io_r_280_b : _GEN_4459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4461 = 9'h119 == r_count_10_io_out ? io_r_281_b : _GEN_4460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4462 = 9'h11a == r_count_10_io_out ? io_r_282_b : _GEN_4461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4463 = 9'h11b == r_count_10_io_out ? io_r_283_b : _GEN_4462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4464 = 9'h11c == r_count_10_io_out ? io_r_284_b : _GEN_4463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4465 = 9'h11d == r_count_10_io_out ? io_r_285_b : _GEN_4464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4466 = 9'h11e == r_count_10_io_out ? io_r_286_b : _GEN_4465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4467 = 9'h11f == r_count_10_io_out ? io_r_287_b : _GEN_4466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4468 = 9'h120 == r_count_10_io_out ? io_r_288_b : _GEN_4467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4469 = 9'h121 == r_count_10_io_out ? io_r_289_b : _GEN_4468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4470 = 9'h122 == r_count_10_io_out ? io_r_290_b : _GEN_4469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4471 = 9'h123 == r_count_10_io_out ? io_r_291_b : _GEN_4470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4472 = 9'h124 == r_count_10_io_out ? io_r_292_b : _GEN_4471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4473 = 9'h125 == r_count_10_io_out ? io_r_293_b : _GEN_4472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4474 = 9'h126 == r_count_10_io_out ? io_r_294_b : _GEN_4473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4475 = 9'h127 == r_count_10_io_out ? io_r_295_b : _GEN_4474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4476 = 9'h128 == r_count_10_io_out ? io_r_296_b : _GEN_4475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4477 = 9'h129 == r_count_10_io_out ? io_r_297_b : _GEN_4476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4478 = 9'h12a == r_count_10_io_out ? io_r_298_b : _GEN_4477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4479 = 9'h12b == r_count_10_io_out ? io_r_299_b : _GEN_4478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4480 = 9'h12c == r_count_10_io_out ? io_r_300_b : _GEN_4479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4481 = 9'h12d == r_count_10_io_out ? io_r_301_b : _GEN_4480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4482 = 9'h12e == r_count_10_io_out ? io_r_302_b : _GEN_4481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4483 = 9'h12f == r_count_10_io_out ? io_r_303_b : _GEN_4482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4484 = 9'h130 == r_count_10_io_out ? io_r_304_b : _GEN_4483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4485 = 9'h131 == r_count_10_io_out ? io_r_305_b : _GEN_4484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4486 = 9'h132 == r_count_10_io_out ? io_r_306_b : _GEN_4485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4487 = 9'h133 == r_count_10_io_out ? io_r_307_b : _GEN_4486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4488 = 9'h134 == r_count_10_io_out ? io_r_308_b : _GEN_4487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4489 = 9'h135 == r_count_10_io_out ? io_r_309_b : _GEN_4488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4490 = 9'h136 == r_count_10_io_out ? io_r_310_b : _GEN_4489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4491 = 9'h137 == r_count_10_io_out ? io_r_311_b : _GEN_4490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4492 = 9'h138 == r_count_10_io_out ? io_r_312_b : _GEN_4491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4493 = 9'h139 == r_count_10_io_out ? io_r_313_b : _GEN_4492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4494 = 9'h13a == r_count_10_io_out ? io_r_314_b : _GEN_4493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4495 = 9'h13b == r_count_10_io_out ? io_r_315_b : _GEN_4494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4496 = 9'h13c == r_count_10_io_out ? io_r_316_b : _GEN_4495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4497 = 9'h13d == r_count_10_io_out ? io_r_317_b : _GEN_4496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4498 = 9'h13e == r_count_10_io_out ? io_r_318_b : _GEN_4497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4499 = 9'h13f == r_count_10_io_out ? io_r_319_b : _GEN_4498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4500 = 9'h140 == r_count_10_io_out ? io_r_320_b : _GEN_4499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4501 = 9'h141 == r_count_10_io_out ? io_r_321_b : _GEN_4500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4502 = 9'h142 == r_count_10_io_out ? io_r_322_b : _GEN_4501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4503 = 9'h143 == r_count_10_io_out ? io_r_323_b : _GEN_4502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4504 = 9'h144 == r_count_10_io_out ? io_r_324_b : _GEN_4503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4505 = 9'h145 == r_count_10_io_out ? io_r_325_b : _GEN_4504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4506 = 9'h146 == r_count_10_io_out ? io_r_326_b : _GEN_4505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4507 = 9'h147 == r_count_10_io_out ? io_r_327_b : _GEN_4506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4508 = 9'h148 == r_count_10_io_out ? io_r_328_b : _GEN_4507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4509 = 9'h149 == r_count_10_io_out ? io_r_329_b : _GEN_4508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4510 = 9'h14a == r_count_10_io_out ? io_r_330_b : _GEN_4509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4511 = 9'h14b == r_count_10_io_out ? io_r_331_b : _GEN_4510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4512 = 9'h14c == r_count_10_io_out ? io_r_332_b : _GEN_4511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4513 = 9'h14d == r_count_10_io_out ? io_r_333_b : _GEN_4512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4514 = 9'h14e == r_count_10_io_out ? io_r_334_b : _GEN_4513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4515 = 9'h14f == r_count_10_io_out ? io_r_335_b : _GEN_4514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4516 = 9'h150 == r_count_10_io_out ? io_r_336_b : _GEN_4515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4517 = 9'h151 == r_count_10_io_out ? io_r_337_b : _GEN_4516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4518 = 9'h152 == r_count_10_io_out ? io_r_338_b : _GEN_4517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4519 = 9'h153 == r_count_10_io_out ? io_r_339_b : _GEN_4518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4520 = 9'h154 == r_count_10_io_out ? io_r_340_b : _GEN_4519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4521 = 9'h155 == r_count_10_io_out ? io_r_341_b : _GEN_4520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4522 = 9'h156 == r_count_10_io_out ? io_r_342_b : _GEN_4521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4523 = 9'h157 == r_count_10_io_out ? io_r_343_b : _GEN_4522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4524 = 9'h158 == r_count_10_io_out ? io_r_344_b : _GEN_4523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4525 = 9'h159 == r_count_10_io_out ? io_r_345_b : _GEN_4524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4526 = 9'h15a == r_count_10_io_out ? io_r_346_b : _GEN_4525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4527 = 9'h15b == r_count_10_io_out ? io_r_347_b : _GEN_4526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4528 = 9'h15c == r_count_10_io_out ? io_r_348_b : _GEN_4527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4529 = 9'h15d == r_count_10_io_out ? io_r_349_b : _GEN_4528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4530 = 9'h15e == r_count_10_io_out ? io_r_350_b : _GEN_4529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4531 = 9'h15f == r_count_10_io_out ? io_r_351_b : _GEN_4530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4532 = 9'h160 == r_count_10_io_out ? io_r_352_b : _GEN_4531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4533 = 9'h161 == r_count_10_io_out ? io_r_353_b : _GEN_4532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4534 = 9'h162 == r_count_10_io_out ? io_r_354_b : _GEN_4533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4535 = 9'h163 == r_count_10_io_out ? io_r_355_b : _GEN_4534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4536 = 9'h164 == r_count_10_io_out ? io_r_356_b : _GEN_4535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4537 = 9'h165 == r_count_10_io_out ? io_r_357_b : _GEN_4536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4538 = 9'h166 == r_count_10_io_out ? io_r_358_b : _GEN_4537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4539 = 9'h167 == r_count_10_io_out ? io_r_359_b : _GEN_4538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4540 = 9'h168 == r_count_10_io_out ? io_r_360_b : _GEN_4539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4541 = 9'h169 == r_count_10_io_out ? io_r_361_b : _GEN_4540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4542 = 9'h16a == r_count_10_io_out ? io_r_362_b : _GEN_4541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4543 = 9'h16b == r_count_10_io_out ? io_r_363_b : _GEN_4542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4544 = 9'h16c == r_count_10_io_out ? io_r_364_b : _GEN_4543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4545 = 9'h16d == r_count_10_io_out ? io_r_365_b : _GEN_4544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4546 = 9'h16e == r_count_10_io_out ? io_r_366_b : _GEN_4545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4547 = 9'h16f == r_count_10_io_out ? io_r_367_b : _GEN_4546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4548 = 9'h170 == r_count_10_io_out ? io_r_368_b : _GEN_4547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4549 = 9'h171 == r_count_10_io_out ? io_r_369_b : _GEN_4548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4550 = 9'h172 == r_count_10_io_out ? io_r_370_b : _GEN_4549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4551 = 9'h173 == r_count_10_io_out ? io_r_371_b : _GEN_4550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4552 = 9'h174 == r_count_10_io_out ? io_r_372_b : _GEN_4551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4553 = 9'h175 == r_count_10_io_out ? io_r_373_b : _GEN_4552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4554 = 9'h176 == r_count_10_io_out ? io_r_374_b : _GEN_4553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4555 = 9'h177 == r_count_10_io_out ? io_r_375_b : _GEN_4554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4556 = 9'h178 == r_count_10_io_out ? io_r_376_b : _GEN_4555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4557 = 9'h179 == r_count_10_io_out ? io_r_377_b : _GEN_4556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4558 = 9'h17a == r_count_10_io_out ? io_r_378_b : _GEN_4557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4559 = 9'h17b == r_count_10_io_out ? io_r_379_b : _GEN_4558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4560 = 9'h17c == r_count_10_io_out ? io_r_380_b : _GEN_4559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4561 = 9'h17d == r_count_10_io_out ? io_r_381_b : _GEN_4560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4562 = 9'h17e == r_count_10_io_out ? io_r_382_b : _GEN_4561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4563 = 9'h17f == r_count_10_io_out ? io_r_383_b : _GEN_4562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4564 = 9'h180 == r_count_10_io_out ? io_r_384_b : _GEN_4563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4565 = 9'h181 == r_count_10_io_out ? io_r_385_b : _GEN_4564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4566 = 9'h182 == r_count_10_io_out ? io_r_386_b : _GEN_4565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4567 = 9'h183 == r_count_10_io_out ? io_r_387_b : _GEN_4566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4568 = 9'h184 == r_count_10_io_out ? io_r_388_b : _GEN_4567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4569 = 9'h185 == r_count_10_io_out ? io_r_389_b : _GEN_4568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4570 = 9'h186 == r_count_10_io_out ? io_r_390_b : _GEN_4569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4571 = 9'h187 == r_count_10_io_out ? io_r_391_b : _GEN_4570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4572 = 9'h188 == r_count_10_io_out ? io_r_392_b : _GEN_4571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4573 = 9'h189 == r_count_10_io_out ? io_r_393_b : _GEN_4572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4574 = 9'h18a == r_count_10_io_out ? io_r_394_b : _GEN_4573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4575 = 9'h18b == r_count_10_io_out ? io_r_395_b : _GEN_4574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4576 = 9'h18c == r_count_10_io_out ? io_r_396_b : _GEN_4575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4577 = 9'h18d == r_count_10_io_out ? io_r_397_b : _GEN_4576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4578 = 9'h18e == r_count_10_io_out ? io_r_398_b : _GEN_4577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4581 = 9'h1 == r_count_11_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4582 = 9'h2 == r_count_11_io_out ? io_r_2_b : _GEN_4581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4583 = 9'h3 == r_count_11_io_out ? io_r_3_b : _GEN_4582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4584 = 9'h4 == r_count_11_io_out ? io_r_4_b : _GEN_4583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4585 = 9'h5 == r_count_11_io_out ? io_r_5_b : _GEN_4584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4586 = 9'h6 == r_count_11_io_out ? io_r_6_b : _GEN_4585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4587 = 9'h7 == r_count_11_io_out ? io_r_7_b : _GEN_4586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4588 = 9'h8 == r_count_11_io_out ? io_r_8_b : _GEN_4587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4589 = 9'h9 == r_count_11_io_out ? io_r_9_b : _GEN_4588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4590 = 9'ha == r_count_11_io_out ? io_r_10_b : _GEN_4589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4591 = 9'hb == r_count_11_io_out ? io_r_11_b : _GEN_4590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4592 = 9'hc == r_count_11_io_out ? io_r_12_b : _GEN_4591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4593 = 9'hd == r_count_11_io_out ? io_r_13_b : _GEN_4592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4594 = 9'he == r_count_11_io_out ? io_r_14_b : _GEN_4593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4595 = 9'hf == r_count_11_io_out ? io_r_15_b : _GEN_4594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4596 = 9'h10 == r_count_11_io_out ? io_r_16_b : _GEN_4595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4597 = 9'h11 == r_count_11_io_out ? io_r_17_b : _GEN_4596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4598 = 9'h12 == r_count_11_io_out ? io_r_18_b : _GEN_4597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4599 = 9'h13 == r_count_11_io_out ? io_r_19_b : _GEN_4598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4600 = 9'h14 == r_count_11_io_out ? io_r_20_b : _GEN_4599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4601 = 9'h15 == r_count_11_io_out ? io_r_21_b : _GEN_4600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4602 = 9'h16 == r_count_11_io_out ? io_r_22_b : _GEN_4601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4603 = 9'h17 == r_count_11_io_out ? io_r_23_b : _GEN_4602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4604 = 9'h18 == r_count_11_io_out ? io_r_24_b : _GEN_4603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4605 = 9'h19 == r_count_11_io_out ? io_r_25_b : _GEN_4604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4606 = 9'h1a == r_count_11_io_out ? io_r_26_b : _GEN_4605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4607 = 9'h1b == r_count_11_io_out ? io_r_27_b : _GEN_4606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4608 = 9'h1c == r_count_11_io_out ? io_r_28_b : _GEN_4607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4609 = 9'h1d == r_count_11_io_out ? io_r_29_b : _GEN_4608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4610 = 9'h1e == r_count_11_io_out ? io_r_30_b : _GEN_4609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4611 = 9'h1f == r_count_11_io_out ? io_r_31_b : _GEN_4610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4612 = 9'h20 == r_count_11_io_out ? io_r_32_b : _GEN_4611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4613 = 9'h21 == r_count_11_io_out ? io_r_33_b : _GEN_4612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4614 = 9'h22 == r_count_11_io_out ? io_r_34_b : _GEN_4613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4615 = 9'h23 == r_count_11_io_out ? io_r_35_b : _GEN_4614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4616 = 9'h24 == r_count_11_io_out ? io_r_36_b : _GEN_4615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4617 = 9'h25 == r_count_11_io_out ? io_r_37_b : _GEN_4616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4618 = 9'h26 == r_count_11_io_out ? io_r_38_b : _GEN_4617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4619 = 9'h27 == r_count_11_io_out ? io_r_39_b : _GEN_4618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4620 = 9'h28 == r_count_11_io_out ? io_r_40_b : _GEN_4619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4621 = 9'h29 == r_count_11_io_out ? io_r_41_b : _GEN_4620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4622 = 9'h2a == r_count_11_io_out ? io_r_42_b : _GEN_4621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4623 = 9'h2b == r_count_11_io_out ? io_r_43_b : _GEN_4622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4624 = 9'h2c == r_count_11_io_out ? io_r_44_b : _GEN_4623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4625 = 9'h2d == r_count_11_io_out ? io_r_45_b : _GEN_4624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4626 = 9'h2e == r_count_11_io_out ? io_r_46_b : _GEN_4625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4627 = 9'h2f == r_count_11_io_out ? io_r_47_b : _GEN_4626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4628 = 9'h30 == r_count_11_io_out ? io_r_48_b : _GEN_4627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4629 = 9'h31 == r_count_11_io_out ? io_r_49_b : _GEN_4628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4630 = 9'h32 == r_count_11_io_out ? io_r_50_b : _GEN_4629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4631 = 9'h33 == r_count_11_io_out ? io_r_51_b : _GEN_4630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4632 = 9'h34 == r_count_11_io_out ? io_r_52_b : _GEN_4631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4633 = 9'h35 == r_count_11_io_out ? io_r_53_b : _GEN_4632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4634 = 9'h36 == r_count_11_io_out ? io_r_54_b : _GEN_4633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4635 = 9'h37 == r_count_11_io_out ? io_r_55_b : _GEN_4634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4636 = 9'h38 == r_count_11_io_out ? io_r_56_b : _GEN_4635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4637 = 9'h39 == r_count_11_io_out ? io_r_57_b : _GEN_4636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4638 = 9'h3a == r_count_11_io_out ? io_r_58_b : _GEN_4637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4639 = 9'h3b == r_count_11_io_out ? io_r_59_b : _GEN_4638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4640 = 9'h3c == r_count_11_io_out ? io_r_60_b : _GEN_4639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4641 = 9'h3d == r_count_11_io_out ? io_r_61_b : _GEN_4640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4642 = 9'h3e == r_count_11_io_out ? io_r_62_b : _GEN_4641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4643 = 9'h3f == r_count_11_io_out ? io_r_63_b : _GEN_4642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4644 = 9'h40 == r_count_11_io_out ? io_r_64_b : _GEN_4643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4645 = 9'h41 == r_count_11_io_out ? io_r_65_b : _GEN_4644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4646 = 9'h42 == r_count_11_io_out ? io_r_66_b : _GEN_4645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4647 = 9'h43 == r_count_11_io_out ? io_r_67_b : _GEN_4646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4648 = 9'h44 == r_count_11_io_out ? io_r_68_b : _GEN_4647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4649 = 9'h45 == r_count_11_io_out ? io_r_69_b : _GEN_4648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4650 = 9'h46 == r_count_11_io_out ? io_r_70_b : _GEN_4649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4651 = 9'h47 == r_count_11_io_out ? io_r_71_b : _GEN_4650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4652 = 9'h48 == r_count_11_io_out ? io_r_72_b : _GEN_4651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4653 = 9'h49 == r_count_11_io_out ? io_r_73_b : _GEN_4652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4654 = 9'h4a == r_count_11_io_out ? io_r_74_b : _GEN_4653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4655 = 9'h4b == r_count_11_io_out ? io_r_75_b : _GEN_4654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4656 = 9'h4c == r_count_11_io_out ? io_r_76_b : _GEN_4655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4657 = 9'h4d == r_count_11_io_out ? io_r_77_b : _GEN_4656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4658 = 9'h4e == r_count_11_io_out ? io_r_78_b : _GEN_4657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4659 = 9'h4f == r_count_11_io_out ? io_r_79_b : _GEN_4658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4660 = 9'h50 == r_count_11_io_out ? io_r_80_b : _GEN_4659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4661 = 9'h51 == r_count_11_io_out ? io_r_81_b : _GEN_4660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4662 = 9'h52 == r_count_11_io_out ? io_r_82_b : _GEN_4661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4663 = 9'h53 == r_count_11_io_out ? io_r_83_b : _GEN_4662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4664 = 9'h54 == r_count_11_io_out ? io_r_84_b : _GEN_4663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4665 = 9'h55 == r_count_11_io_out ? io_r_85_b : _GEN_4664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4666 = 9'h56 == r_count_11_io_out ? io_r_86_b : _GEN_4665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4667 = 9'h57 == r_count_11_io_out ? io_r_87_b : _GEN_4666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4668 = 9'h58 == r_count_11_io_out ? io_r_88_b : _GEN_4667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4669 = 9'h59 == r_count_11_io_out ? io_r_89_b : _GEN_4668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4670 = 9'h5a == r_count_11_io_out ? io_r_90_b : _GEN_4669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4671 = 9'h5b == r_count_11_io_out ? io_r_91_b : _GEN_4670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4672 = 9'h5c == r_count_11_io_out ? io_r_92_b : _GEN_4671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4673 = 9'h5d == r_count_11_io_out ? io_r_93_b : _GEN_4672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4674 = 9'h5e == r_count_11_io_out ? io_r_94_b : _GEN_4673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4675 = 9'h5f == r_count_11_io_out ? io_r_95_b : _GEN_4674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4676 = 9'h60 == r_count_11_io_out ? io_r_96_b : _GEN_4675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4677 = 9'h61 == r_count_11_io_out ? io_r_97_b : _GEN_4676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4678 = 9'h62 == r_count_11_io_out ? io_r_98_b : _GEN_4677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4679 = 9'h63 == r_count_11_io_out ? io_r_99_b : _GEN_4678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4680 = 9'h64 == r_count_11_io_out ? io_r_100_b : _GEN_4679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4681 = 9'h65 == r_count_11_io_out ? io_r_101_b : _GEN_4680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4682 = 9'h66 == r_count_11_io_out ? io_r_102_b : _GEN_4681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4683 = 9'h67 == r_count_11_io_out ? io_r_103_b : _GEN_4682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4684 = 9'h68 == r_count_11_io_out ? io_r_104_b : _GEN_4683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4685 = 9'h69 == r_count_11_io_out ? io_r_105_b : _GEN_4684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4686 = 9'h6a == r_count_11_io_out ? io_r_106_b : _GEN_4685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4687 = 9'h6b == r_count_11_io_out ? io_r_107_b : _GEN_4686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4688 = 9'h6c == r_count_11_io_out ? io_r_108_b : _GEN_4687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4689 = 9'h6d == r_count_11_io_out ? io_r_109_b : _GEN_4688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4690 = 9'h6e == r_count_11_io_out ? io_r_110_b : _GEN_4689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4691 = 9'h6f == r_count_11_io_out ? io_r_111_b : _GEN_4690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4692 = 9'h70 == r_count_11_io_out ? io_r_112_b : _GEN_4691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4693 = 9'h71 == r_count_11_io_out ? io_r_113_b : _GEN_4692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4694 = 9'h72 == r_count_11_io_out ? io_r_114_b : _GEN_4693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4695 = 9'h73 == r_count_11_io_out ? io_r_115_b : _GEN_4694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4696 = 9'h74 == r_count_11_io_out ? io_r_116_b : _GEN_4695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4697 = 9'h75 == r_count_11_io_out ? io_r_117_b : _GEN_4696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4698 = 9'h76 == r_count_11_io_out ? io_r_118_b : _GEN_4697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4699 = 9'h77 == r_count_11_io_out ? io_r_119_b : _GEN_4698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4700 = 9'h78 == r_count_11_io_out ? io_r_120_b : _GEN_4699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4701 = 9'h79 == r_count_11_io_out ? io_r_121_b : _GEN_4700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4702 = 9'h7a == r_count_11_io_out ? io_r_122_b : _GEN_4701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4703 = 9'h7b == r_count_11_io_out ? io_r_123_b : _GEN_4702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4704 = 9'h7c == r_count_11_io_out ? io_r_124_b : _GEN_4703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4705 = 9'h7d == r_count_11_io_out ? io_r_125_b : _GEN_4704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4706 = 9'h7e == r_count_11_io_out ? io_r_126_b : _GEN_4705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4707 = 9'h7f == r_count_11_io_out ? io_r_127_b : _GEN_4706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4708 = 9'h80 == r_count_11_io_out ? io_r_128_b : _GEN_4707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4709 = 9'h81 == r_count_11_io_out ? io_r_129_b : _GEN_4708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4710 = 9'h82 == r_count_11_io_out ? io_r_130_b : _GEN_4709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4711 = 9'h83 == r_count_11_io_out ? io_r_131_b : _GEN_4710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4712 = 9'h84 == r_count_11_io_out ? io_r_132_b : _GEN_4711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4713 = 9'h85 == r_count_11_io_out ? io_r_133_b : _GEN_4712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4714 = 9'h86 == r_count_11_io_out ? io_r_134_b : _GEN_4713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4715 = 9'h87 == r_count_11_io_out ? io_r_135_b : _GEN_4714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4716 = 9'h88 == r_count_11_io_out ? io_r_136_b : _GEN_4715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4717 = 9'h89 == r_count_11_io_out ? io_r_137_b : _GEN_4716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4718 = 9'h8a == r_count_11_io_out ? io_r_138_b : _GEN_4717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4719 = 9'h8b == r_count_11_io_out ? io_r_139_b : _GEN_4718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4720 = 9'h8c == r_count_11_io_out ? io_r_140_b : _GEN_4719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4721 = 9'h8d == r_count_11_io_out ? io_r_141_b : _GEN_4720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4722 = 9'h8e == r_count_11_io_out ? io_r_142_b : _GEN_4721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4723 = 9'h8f == r_count_11_io_out ? io_r_143_b : _GEN_4722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4724 = 9'h90 == r_count_11_io_out ? io_r_144_b : _GEN_4723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4725 = 9'h91 == r_count_11_io_out ? io_r_145_b : _GEN_4724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4726 = 9'h92 == r_count_11_io_out ? io_r_146_b : _GEN_4725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4727 = 9'h93 == r_count_11_io_out ? io_r_147_b : _GEN_4726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4728 = 9'h94 == r_count_11_io_out ? io_r_148_b : _GEN_4727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4729 = 9'h95 == r_count_11_io_out ? io_r_149_b : _GEN_4728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4730 = 9'h96 == r_count_11_io_out ? io_r_150_b : _GEN_4729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4731 = 9'h97 == r_count_11_io_out ? io_r_151_b : _GEN_4730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4732 = 9'h98 == r_count_11_io_out ? io_r_152_b : _GEN_4731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4733 = 9'h99 == r_count_11_io_out ? io_r_153_b : _GEN_4732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4734 = 9'h9a == r_count_11_io_out ? io_r_154_b : _GEN_4733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4735 = 9'h9b == r_count_11_io_out ? io_r_155_b : _GEN_4734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4736 = 9'h9c == r_count_11_io_out ? io_r_156_b : _GEN_4735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4737 = 9'h9d == r_count_11_io_out ? io_r_157_b : _GEN_4736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4738 = 9'h9e == r_count_11_io_out ? io_r_158_b : _GEN_4737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4739 = 9'h9f == r_count_11_io_out ? io_r_159_b : _GEN_4738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4740 = 9'ha0 == r_count_11_io_out ? io_r_160_b : _GEN_4739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4741 = 9'ha1 == r_count_11_io_out ? io_r_161_b : _GEN_4740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4742 = 9'ha2 == r_count_11_io_out ? io_r_162_b : _GEN_4741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4743 = 9'ha3 == r_count_11_io_out ? io_r_163_b : _GEN_4742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4744 = 9'ha4 == r_count_11_io_out ? io_r_164_b : _GEN_4743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4745 = 9'ha5 == r_count_11_io_out ? io_r_165_b : _GEN_4744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4746 = 9'ha6 == r_count_11_io_out ? io_r_166_b : _GEN_4745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4747 = 9'ha7 == r_count_11_io_out ? io_r_167_b : _GEN_4746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4748 = 9'ha8 == r_count_11_io_out ? io_r_168_b : _GEN_4747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4749 = 9'ha9 == r_count_11_io_out ? io_r_169_b : _GEN_4748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4750 = 9'haa == r_count_11_io_out ? io_r_170_b : _GEN_4749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4751 = 9'hab == r_count_11_io_out ? io_r_171_b : _GEN_4750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4752 = 9'hac == r_count_11_io_out ? io_r_172_b : _GEN_4751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4753 = 9'had == r_count_11_io_out ? io_r_173_b : _GEN_4752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4754 = 9'hae == r_count_11_io_out ? io_r_174_b : _GEN_4753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4755 = 9'haf == r_count_11_io_out ? io_r_175_b : _GEN_4754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4756 = 9'hb0 == r_count_11_io_out ? io_r_176_b : _GEN_4755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4757 = 9'hb1 == r_count_11_io_out ? io_r_177_b : _GEN_4756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4758 = 9'hb2 == r_count_11_io_out ? io_r_178_b : _GEN_4757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4759 = 9'hb3 == r_count_11_io_out ? io_r_179_b : _GEN_4758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4760 = 9'hb4 == r_count_11_io_out ? io_r_180_b : _GEN_4759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4761 = 9'hb5 == r_count_11_io_out ? io_r_181_b : _GEN_4760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4762 = 9'hb6 == r_count_11_io_out ? io_r_182_b : _GEN_4761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4763 = 9'hb7 == r_count_11_io_out ? io_r_183_b : _GEN_4762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4764 = 9'hb8 == r_count_11_io_out ? io_r_184_b : _GEN_4763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4765 = 9'hb9 == r_count_11_io_out ? io_r_185_b : _GEN_4764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4766 = 9'hba == r_count_11_io_out ? io_r_186_b : _GEN_4765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4767 = 9'hbb == r_count_11_io_out ? io_r_187_b : _GEN_4766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4768 = 9'hbc == r_count_11_io_out ? io_r_188_b : _GEN_4767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4769 = 9'hbd == r_count_11_io_out ? io_r_189_b : _GEN_4768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4770 = 9'hbe == r_count_11_io_out ? io_r_190_b : _GEN_4769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4771 = 9'hbf == r_count_11_io_out ? io_r_191_b : _GEN_4770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4772 = 9'hc0 == r_count_11_io_out ? io_r_192_b : _GEN_4771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4773 = 9'hc1 == r_count_11_io_out ? io_r_193_b : _GEN_4772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4774 = 9'hc2 == r_count_11_io_out ? io_r_194_b : _GEN_4773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4775 = 9'hc3 == r_count_11_io_out ? io_r_195_b : _GEN_4774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4776 = 9'hc4 == r_count_11_io_out ? io_r_196_b : _GEN_4775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4777 = 9'hc5 == r_count_11_io_out ? io_r_197_b : _GEN_4776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4778 = 9'hc6 == r_count_11_io_out ? io_r_198_b : _GEN_4777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4779 = 9'hc7 == r_count_11_io_out ? io_r_199_b : _GEN_4778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4780 = 9'hc8 == r_count_11_io_out ? io_r_200_b : _GEN_4779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4781 = 9'hc9 == r_count_11_io_out ? io_r_201_b : _GEN_4780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4782 = 9'hca == r_count_11_io_out ? io_r_202_b : _GEN_4781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4783 = 9'hcb == r_count_11_io_out ? io_r_203_b : _GEN_4782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4784 = 9'hcc == r_count_11_io_out ? io_r_204_b : _GEN_4783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4785 = 9'hcd == r_count_11_io_out ? io_r_205_b : _GEN_4784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4786 = 9'hce == r_count_11_io_out ? io_r_206_b : _GEN_4785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4787 = 9'hcf == r_count_11_io_out ? io_r_207_b : _GEN_4786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4788 = 9'hd0 == r_count_11_io_out ? io_r_208_b : _GEN_4787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4789 = 9'hd1 == r_count_11_io_out ? io_r_209_b : _GEN_4788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4790 = 9'hd2 == r_count_11_io_out ? io_r_210_b : _GEN_4789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4791 = 9'hd3 == r_count_11_io_out ? io_r_211_b : _GEN_4790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4792 = 9'hd4 == r_count_11_io_out ? io_r_212_b : _GEN_4791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4793 = 9'hd5 == r_count_11_io_out ? io_r_213_b : _GEN_4792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4794 = 9'hd6 == r_count_11_io_out ? io_r_214_b : _GEN_4793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4795 = 9'hd7 == r_count_11_io_out ? io_r_215_b : _GEN_4794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4796 = 9'hd8 == r_count_11_io_out ? io_r_216_b : _GEN_4795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4797 = 9'hd9 == r_count_11_io_out ? io_r_217_b : _GEN_4796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4798 = 9'hda == r_count_11_io_out ? io_r_218_b : _GEN_4797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4799 = 9'hdb == r_count_11_io_out ? io_r_219_b : _GEN_4798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4800 = 9'hdc == r_count_11_io_out ? io_r_220_b : _GEN_4799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4801 = 9'hdd == r_count_11_io_out ? io_r_221_b : _GEN_4800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4802 = 9'hde == r_count_11_io_out ? io_r_222_b : _GEN_4801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4803 = 9'hdf == r_count_11_io_out ? io_r_223_b : _GEN_4802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4804 = 9'he0 == r_count_11_io_out ? io_r_224_b : _GEN_4803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4805 = 9'he1 == r_count_11_io_out ? io_r_225_b : _GEN_4804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4806 = 9'he2 == r_count_11_io_out ? io_r_226_b : _GEN_4805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4807 = 9'he3 == r_count_11_io_out ? io_r_227_b : _GEN_4806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4808 = 9'he4 == r_count_11_io_out ? io_r_228_b : _GEN_4807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4809 = 9'he5 == r_count_11_io_out ? io_r_229_b : _GEN_4808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4810 = 9'he6 == r_count_11_io_out ? io_r_230_b : _GEN_4809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4811 = 9'he7 == r_count_11_io_out ? io_r_231_b : _GEN_4810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4812 = 9'he8 == r_count_11_io_out ? io_r_232_b : _GEN_4811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4813 = 9'he9 == r_count_11_io_out ? io_r_233_b : _GEN_4812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4814 = 9'hea == r_count_11_io_out ? io_r_234_b : _GEN_4813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4815 = 9'heb == r_count_11_io_out ? io_r_235_b : _GEN_4814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4816 = 9'hec == r_count_11_io_out ? io_r_236_b : _GEN_4815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4817 = 9'hed == r_count_11_io_out ? io_r_237_b : _GEN_4816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4818 = 9'hee == r_count_11_io_out ? io_r_238_b : _GEN_4817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4819 = 9'hef == r_count_11_io_out ? io_r_239_b : _GEN_4818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4820 = 9'hf0 == r_count_11_io_out ? io_r_240_b : _GEN_4819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4821 = 9'hf1 == r_count_11_io_out ? io_r_241_b : _GEN_4820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4822 = 9'hf2 == r_count_11_io_out ? io_r_242_b : _GEN_4821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4823 = 9'hf3 == r_count_11_io_out ? io_r_243_b : _GEN_4822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4824 = 9'hf4 == r_count_11_io_out ? io_r_244_b : _GEN_4823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4825 = 9'hf5 == r_count_11_io_out ? io_r_245_b : _GEN_4824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4826 = 9'hf6 == r_count_11_io_out ? io_r_246_b : _GEN_4825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4827 = 9'hf7 == r_count_11_io_out ? io_r_247_b : _GEN_4826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4828 = 9'hf8 == r_count_11_io_out ? io_r_248_b : _GEN_4827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4829 = 9'hf9 == r_count_11_io_out ? io_r_249_b : _GEN_4828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4830 = 9'hfa == r_count_11_io_out ? io_r_250_b : _GEN_4829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4831 = 9'hfb == r_count_11_io_out ? io_r_251_b : _GEN_4830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4832 = 9'hfc == r_count_11_io_out ? io_r_252_b : _GEN_4831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4833 = 9'hfd == r_count_11_io_out ? io_r_253_b : _GEN_4832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4834 = 9'hfe == r_count_11_io_out ? io_r_254_b : _GEN_4833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4835 = 9'hff == r_count_11_io_out ? io_r_255_b : _GEN_4834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4836 = 9'h100 == r_count_11_io_out ? io_r_256_b : _GEN_4835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4837 = 9'h101 == r_count_11_io_out ? io_r_257_b : _GEN_4836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4838 = 9'h102 == r_count_11_io_out ? io_r_258_b : _GEN_4837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4839 = 9'h103 == r_count_11_io_out ? io_r_259_b : _GEN_4838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4840 = 9'h104 == r_count_11_io_out ? io_r_260_b : _GEN_4839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4841 = 9'h105 == r_count_11_io_out ? io_r_261_b : _GEN_4840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4842 = 9'h106 == r_count_11_io_out ? io_r_262_b : _GEN_4841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4843 = 9'h107 == r_count_11_io_out ? io_r_263_b : _GEN_4842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4844 = 9'h108 == r_count_11_io_out ? io_r_264_b : _GEN_4843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4845 = 9'h109 == r_count_11_io_out ? io_r_265_b : _GEN_4844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4846 = 9'h10a == r_count_11_io_out ? io_r_266_b : _GEN_4845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4847 = 9'h10b == r_count_11_io_out ? io_r_267_b : _GEN_4846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4848 = 9'h10c == r_count_11_io_out ? io_r_268_b : _GEN_4847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4849 = 9'h10d == r_count_11_io_out ? io_r_269_b : _GEN_4848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4850 = 9'h10e == r_count_11_io_out ? io_r_270_b : _GEN_4849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4851 = 9'h10f == r_count_11_io_out ? io_r_271_b : _GEN_4850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4852 = 9'h110 == r_count_11_io_out ? io_r_272_b : _GEN_4851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4853 = 9'h111 == r_count_11_io_out ? io_r_273_b : _GEN_4852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4854 = 9'h112 == r_count_11_io_out ? io_r_274_b : _GEN_4853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4855 = 9'h113 == r_count_11_io_out ? io_r_275_b : _GEN_4854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4856 = 9'h114 == r_count_11_io_out ? io_r_276_b : _GEN_4855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4857 = 9'h115 == r_count_11_io_out ? io_r_277_b : _GEN_4856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4858 = 9'h116 == r_count_11_io_out ? io_r_278_b : _GEN_4857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4859 = 9'h117 == r_count_11_io_out ? io_r_279_b : _GEN_4858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4860 = 9'h118 == r_count_11_io_out ? io_r_280_b : _GEN_4859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4861 = 9'h119 == r_count_11_io_out ? io_r_281_b : _GEN_4860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4862 = 9'h11a == r_count_11_io_out ? io_r_282_b : _GEN_4861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4863 = 9'h11b == r_count_11_io_out ? io_r_283_b : _GEN_4862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4864 = 9'h11c == r_count_11_io_out ? io_r_284_b : _GEN_4863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4865 = 9'h11d == r_count_11_io_out ? io_r_285_b : _GEN_4864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4866 = 9'h11e == r_count_11_io_out ? io_r_286_b : _GEN_4865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4867 = 9'h11f == r_count_11_io_out ? io_r_287_b : _GEN_4866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4868 = 9'h120 == r_count_11_io_out ? io_r_288_b : _GEN_4867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4869 = 9'h121 == r_count_11_io_out ? io_r_289_b : _GEN_4868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4870 = 9'h122 == r_count_11_io_out ? io_r_290_b : _GEN_4869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4871 = 9'h123 == r_count_11_io_out ? io_r_291_b : _GEN_4870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4872 = 9'h124 == r_count_11_io_out ? io_r_292_b : _GEN_4871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4873 = 9'h125 == r_count_11_io_out ? io_r_293_b : _GEN_4872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4874 = 9'h126 == r_count_11_io_out ? io_r_294_b : _GEN_4873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4875 = 9'h127 == r_count_11_io_out ? io_r_295_b : _GEN_4874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4876 = 9'h128 == r_count_11_io_out ? io_r_296_b : _GEN_4875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4877 = 9'h129 == r_count_11_io_out ? io_r_297_b : _GEN_4876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4878 = 9'h12a == r_count_11_io_out ? io_r_298_b : _GEN_4877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4879 = 9'h12b == r_count_11_io_out ? io_r_299_b : _GEN_4878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4880 = 9'h12c == r_count_11_io_out ? io_r_300_b : _GEN_4879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4881 = 9'h12d == r_count_11_io_out ? io_r_301_b : _GEN_4880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4882 = 9'h12e == r_count_11_io_out ? io_r_302_b : _GEN_4881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4883 = 9'h12f == r_count_11_io_out ? io_r_303_b : _GEN_4882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4884 = 9'h130 == r_count_11_io_out ? io_r_304_b : _GEN_4883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4885 = 9'h131 == r_count_11_io_out ? io_r_305_b : _GEN_4884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4886 = 9'h132 == r_count_11_io_out ? io_r_306_b : _GEN_4885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4887 = 9'h133 == r_count_11_io_out ? io_r_307_b : _GEN_4886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4888 = 9'h134 == r_count_11_io_out ? io_r_308_b : _GEN_4887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4889 = 9'h135 == r_count_11_io_out ? io_r_309_b : _GEN_4888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4890 = 9'h136 == r_count_11_io_out ? io_r_310_b : _GEN_4889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4891 = 9'h137 == r_count_11_io_out ? io_r_311_b : _GEN_4890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4892 = 9'h138 == r_count_11_io_out ? io_r_312_b : _GEN_4891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4893 = 9'h139 == r_count_11_io_out ? io_r_313_b : _GEN_4892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4894 = 9'h13a == r_count_11_io_out ? io_r_314_b : _GEN_4893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4895 = 9'h13b == r_count_11_io_out ? io_r_315_b : _GEN_4894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4896 = 9'h13c == r_count_11_io_out ? io_r_316_b : _GEN_4895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4897 = 9'h13d == r_count_11_io_out ? io_r_317_b : _GEN_4896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4898 = 9'h13e == r_count_11_io_out ? io_r_318_b : _GEN_4897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4899 = 9'h13f == r_count_11_io_out ? io_r_319_b : _GEN_4898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4900 = 9'h140 == r_count_11_io_out ? io_r_320_b : _GEN_4899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4901 = 9'h141 == r_count_11_io_out ? io_r_321_b : _GEN_4900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4902 = 9'h142 == r_count_11_io_out ? io_r_322_b : _GEN_4901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4903 = 9'h143 == r_count_11_io_out ? io_r_323_b : _GEN_4902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4904 = 9'h144 == r_count_11_io_out ? io_r_324_b : _GEN_4903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4905 = 9'h145 == r_count_11_io_out ? io_r_325_b : _GEN_4904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4906 = 9'h146 == r_count_11_io_out ? io_r_326_b : _GEN_4905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4907 = 9'h147 == r_count_11_io_out ? io_r_327_b : _GEN_4906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4908 = 9'h148 == r_count_11_io_out ? io_r_328_b : _GEN_4907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4909 = 9'h149 == r_count_11_io_out ? io_r_329_b : _GEN_4908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4910 = 9'h14a == r_count_11_io_out ? io_r_330_b : _GEN_4909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4911 = 9'h14b == r_count_11_io_out ? io_r_331_b : _GEN_4910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4912 = 9'h14c == r_count_11_io_out ? io_r_332_b : _GEN_4911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4913 = 9'h14d == r_count_11_io_out ? io_r_333_b : _GEN_4912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4914 = 9'h14e == r_count_11_io_out ? io_r_334_b : _GEN_4913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4915 = 9'h14f == r_count_11_io_out ? io_r_335_b : _GEN_4914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4916 = 9'h150 == r_count_11_io_out ? io_r_336_b : _GEN_4915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4917 = 9'h151 == r_count_11_io_out ? io_r_337_b : _GEN_4916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4918 = 9'h152 == r_count_11_io_out ? io_r_338_b : _GEN_4917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4919 = 9'h153 == r_count_11_io_out ? io_r_339_b : _GEN_4918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4920 = 9'h154 == r_count_11_io_out ? io_r_340_b : _GEN_4919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4921 = 9'h155 == r_count_11_io_out ? io_r_341_b : _GEN_4920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4922 = 9'h156 == r_count_11_io_out ? io_r_342_b : _GEN_4921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4923 = 9'h157 == r_count_11_io_out ? io_r_343_b : _GEN_4922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4924 = 9'h158 == r_count_11_io_out ? io_r_344_b : _GEN_4923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4925 = 9'h159 == r_count_11_io_out ? io_r_345_b : _GEN_4924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4926 = 9'h15a == r_count_11_io_out ? io_r_346_b : _GEN_4925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4927 = 9'h15b == r_count_11_io_out ? io_r_347_b : _GEN_4926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4928 = 9'h15c == r_count_11_io_out ? io_r_348_b : _GEN_4927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4929 = 9'h15d == r_count_11_io_out ? io_r_349_b : _GEN_4928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4930 = 9'h15e == r_count_11_io_out ? io_r_350_b : _GEN_4929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4931 = 9'h15f == r_count_11_io_out ? io_r_351_b : _GEN_4930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4932 = 9'h160 == r_count_11_io_out ? io_r_352_b : _GEN_4931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4933 = 9'h161 == r_count_11_io_out ? io_r_353_b : _GEN_4932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4934 = 9'h162 == r_count_11_io_out ? io_r_354_b : _GEN_4933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4935 = 9'h163 == r_count_11_io_out ? io_r_355_b : _GEN_4934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4936 = 9'h164 == r_count_11_io_out ? io_r_356_b : _GEN_4935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4937 = 9'h165 == r_count_11_io_out ? io_r_357_b : _GEN_4936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4938 = 9'h166 == r_count_11_io_out ? io_r_358_b : _GEN_4937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4939 = 9'h167 == r_count_11_io_out ? io_r_359_b : _GEN_4938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4940 = 9'h168 == r_count_11_io_out ? io_r_360_b : _GEN_4939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4941 = 9'h169 == r_count_11_io_out ? io_r_361_b : _GEN_4940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4942 = 9'h16a == r_count_11_io_out ? io_r_362_b : _GEN_4941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4943 = 9'h16b == r_count_11_io_out ? io_r_363_b : _GEN_4942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4944 = 9'h16c == r_count_11_io_out ? io_r_364_b : _GEN_4943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4945 = 9'h16d == r_count_11_io_out ? io_r_365_b : _GEN_4944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4946 = 9'h16e == r_count_11_io_out ? io_r_366_b : _GEN_4945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4947 = 9'h16f == r_count_11_io_out ? io_r_367_b : _GEN_4946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4948 = 9'h170 == r_count_11_io_out ? io_r_368_b : _GEN_4947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4949 = 9'h171 == r_count_11_io_out ? io_r_369_b : _GEN_4948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4950 = 9'h172 == r_count_11_io_out ? io_r_370_b : _GEN_4949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4951 = 9'h173 == r_count_11_io_out ? io_r_371_b : _GEN_4950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4952 = 9'h174 == r_count_11_io_out ? io_r_372_b : _GEN_4951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4953 = 9'h175 == r_count_11_io_out ? io_r_373_b : _GEN_4952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4954 = 9'h176 == r_count_11_io_out ? io_r_374_b : _GEN_4953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4955 = 9'h177 == r_count_11_io_out ? io_r_375_b : _GEN_4954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4956 = 9'h178 == r_count_11_io_out ? io_r_376_b : _GEN_4955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4957 = 9'h179 == r_count_11_io_out ? io_r_377_b : _GEN_4956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4958 = 9'h17a == r_count_11_io_out ? io_r_378_b : _GEN_4957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4959 = 9'h17b == r_count_11_io_out ? io_r_379_b : _GEN_4958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4960 = 9'h17c == r_count_11_io_out ? io_r_380_b : _GEN_4959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4961 = 9'h17d == r_count_11_io_out ? io_r_381_b : _GEN_4960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4962 = 9'h17e == r_count_11_io_out ? io_r_382_b : _GEN_4961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4963 = 9'h17f == r_count_11_io_out ? io_r_383_b : _GEN_4962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4964 = 9'h180 == r_count_11_io_out ? io_r_384_b : _GEN_4963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4965 = 9'h181 == r_count_11_io_out ? io_r_385_b : _GEN_4964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4966 = 9'h182 == r_count_11_io_out ? io_r_386_b : _GEN_4965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4967 = 9'h183 == r_count_11_io_out ? io_r_387_b : _GEN_4966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4968 = 9'h184 == r_count_11_io_out ? io_r_388_b : _GEN_4967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4969 = 9'h185 == r_count_11_io_out ? io_r_389_b : _GEN_4968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4970 = 9'h186 == r_count_11_io_out ? io_r_390_b : _GEN_4969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4971 = 9'h187 == r_count_11_io_out ? io_r_391_b : _GEN_4970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4972 = 9'h188 == r_count_11_io_out ? io_r_392_b : _GEN_4971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4973 = 9'h189 == r_count_11_io_out ? io_r_393_b : _GEN_4972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4974 = 9'h18a == r_count_11_io_out ? io_r_394_b : _GEN_4973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4975 = 9'h18b == r_count_11_io_out ? io_r_395_b : _GEN_4974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4976 = 9'h18c == r_count_11_io_out ? io_r_396_b : _GEN_4975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4977 = 9'h18d == r_count_11_io_out ? io_r_397_b : _GEN_4976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4978 = 9'h18e == r_count_11_io_out ? io_r_398_b : _GEN_4977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4981 = 9'h1 == r_count_12_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4982 = 9'h2 == r_count_12_io_out ? io_r_2_b : _GEN_4981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4983 = 9'h3 == r_count_12_io_out ? io_r_3_b : _GEN_4982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4984 = 9'h4 == r_count_12_io_out ? io_r_4_b : _GEN_4983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4985 = 9'h5 == r_count_12_io_out ? io_r_5_b : _GEN_4984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4986 = 9'h6 == r_count_12_io_out ? io_r_6_b : _GEN_4985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4987 = 9'h7 == r_count_12_io_out ? io_r_7_b : _GEN_4986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4988 = 9'h8 == r_count_12_io_out ? io_r_8_b : _GEN_4987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4989 = 9'h9 == r_count_12_io_out ? io_r_9_b : _GEN_4988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4990 = 9'ha == r_count_12_io_out ? io_r_10_b : _GEN_4989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4991 = 9'hb == r_count_12_io_out ? io_r_11_b : _GEN_4990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4992 = 9'hc == r_count_12_io_out ? io_r_12_b : _GEN_4991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4993 = 9'hd == r_count_12_io_out ? io_r_13_b : _GEN_4992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4994 = 9'he == r_count_12_io_out ? io_r_14_b : _GEN_4993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4995 = 9'hf == r_count_12_io_out ? io_r_15_b : _GEN_4994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4996 = 9'h10 == r_count_12_io_out ? io_r_16_b : _GEN_4995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4997 = 9'h11 == r_count_12_io_out ? io_r_17_b : _GEN_4996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4998 = 9'h12 == r_count_12_io_out ? io_r_18_b : _GEN_4997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4999 = 9'h13 == r_count_12_io_out ? io_r_19_b : _GEN_4998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5000 = 9'h14 == r_count_12_io_out ? io_r_20_b : _GEN_4999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5001 = 9'h15 == r_count_12_io_out ? io_r_21_b : _GEN_5000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5002 = 9'h16 == r_count_12_io_out ? io_r_22_b : _GEN_5001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5003 = 9'h17 == r_count_12_io_out ? io_r_23_b : _GEN_5002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5004 = 9'h18 == r_count_12_io_out ? io_r_24_b : _GEN_5003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5005 = 9'h19 == r_count_12_io_out ? io_r_25_b : _GEN_5004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5006 = 9'h1a == r_count_12_io_out ? io_r_26_b : _GEN_5005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5007 = 9'h1b == r_count_12_io_out ? io_r_27_b : _GEN_5006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5008 = 9'h1c == r_count_12_io_out ? io_r_28_b : _GEN_5007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5009 = 9'h1d == r_count_12_io_out ? io_r_29_b : _GEN_5008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5010 = 9'h1e == r_count_12_io_out ? io_r_30_b : _GEN_5009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5011 = 9'h1f == r_count_12_io_out ? io_r_31_b : _GEN_5010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5012 = 9'h20 == r_count_12_io_out ? io_r_32_b : _GEN_5011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5013 = 9'h21 == r_count_12_io_out ? io_r_33_b : _GEN_5012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5014 = 9'h22 == r_count_12_io_out ? io_r_34_b : _GEN_5013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5015 = 9'h23 == r_count_12_io_out ? io_r_35_b : _GEN_5014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5016 = 9'h24 == r_count_12_io_out ? io_r_36_b : _GEN_5015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5017 = 9'h25 == r_count_12_io_out ? io_r_37_b : _GEN_5016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5018 = 9'h26 == r_count_12_io_out ? io_r_38_b : _GEN_5017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5019 = 9'h27 == r_count_12_io_out ? io_r_39_b : _GEN_5018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5020 = 9'h28 == r_count_12_io_out ? io_r_40_b : _GEN_5019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5021 = 9'h29 == r_count_12_io_out ? io_r_41_b : _GEN_5020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5022 = 9'h2a == r_count_12_io_out ? io_r_42_b : _GEN_5021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5023 = 9'h2b == r_count_12_io_out ? io_r_43_b : _GEN_5022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5024 = 9'h2c == r_count_12_io_out ? io_r_44_b : _GEN_5023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5025 = 9'h2d == r_count_12_io_out ? io_r_45_b : _GEN_5024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5026 = 9'h2e == r_count_12_io_out ? io_r_46_b : _GEN_5025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5027 = 9'h2f == r_count_12_io_out ? io_r_47_b : _GEN_5026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5028 = 9'h30 == r_count_12_io_out ? io_r_48_b : _GEN_5027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5029 = 9'h31 == r_count_12_io_out ? io_r_49_b : _GEN_5028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5030 = 9'h32 == r_count_12_io_out ? io_r_50_b : _GEN_5029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5031 = 9'h33 == r_count_12_io_out ? io_r_51_b : _GEN_5030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5032 = 9'h34 == r_count_12_io_out ? io_r_52_b : _GEN_5031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5033 = 9'h35 == r_count_12_io_out ? io_r_53_b : _GEN_5032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5034 = 9'h36 == r_count_12_io_out ? io_r_54_b : _GEN_5033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5035 = 9'h37 == r_count_12_io_out ? io_r_55_b : _GEN_5034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5036 = 9'h38 == r_count_12_io_out ? io_r_56_b : _GEN_5035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5037 = 9'h39 == r_count_12_io_out ? io_r_57_b : _GEN_5036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5038 = 9'h3a == r_count_12_io_out ? io_r_58_b : _GEN_5037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5039 = 9'h3b == r_count_12_io_out ? io_r_59_b : _GEN_5038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5040 = 9'h3c == r_count_12_io_out ? io_r_60_b : _GEN_5039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5041 = 9'h3d == r_count_12_io_out ? io_r_61_b : _GEN_5040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5042 = 9'h3e == r_count_12_io_out ? io_r_62_b : _GEN_5041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5043 = 9'h3f == r_count_12_io_out ? io_r_63_b : _GEN_5042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5044 = 9'h40 == r_count_12_io_out ? io_r_64_b : _GEN_5043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5045 = 9'h41 == r_count_12_io_out ? io_r_65_b : _GEN_5044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5046 = 9'h42 == r_count_12_io_out ? io_r_66_b : _GEN_5045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5047 = 9'h43 == r_count_12_io_out ? io_r_67_b : _GEN_5046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5048 = 9'h44 == r_count_12_io_out ? io_r_68_b : _GEN_5047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5049 = 9'h45 == r_count_12_io_out ? io_r_69_b : _GEN_5048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5050 = 9'h46 == r_count_12_io_out ? io_r_70_b : _GEN_5049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5051 = 9'h47 == r_count_12_io_out ? io_r_71_b : _GEN_5050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5052 = 9'h48 == r_count_12_io_out ? io_r_72_b : _GEN_5051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5053 = 9'h49 == r_count_12_io_out ? io_r_73_b : _GEN_5052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5054 = 9'h4a == r_count_12_io_out ? io_r_74_b : _GEN_5053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5055 = 9'h4b == r_count_12_io_out ? io_r_75_b : _GEN_5054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5056 = 9'h4c == r_count_12_io_out ? io_r_76_b : _GEN_5055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5057 = 9'h4d == r_count_12_io_out ? io_r_77_b : _GEN_5056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5058 = 9'h4e == r_count_12_io_out ? io_r_78_b : _GEN_5057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5059 = 9'h4f == r_count_12_io_out ? io_r_79_b : _GEN_5058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5060 = 9'h50 == r_count_12_io_out ? io_r_80_b : _GEN_5059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5061 = 9'h51 == r_count_12_io_out ? io_r_81_b : _GEN_5060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5062 = 9'h52 == r_count_12_io_out ? io_r_82_b : _GEN_5061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5063 = 9'h53 == r_count_12_io_out ? io_r_83_b : _GEN_5062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5064 = 9'h54 == r_count_12_io_out ? io_r_84_b : _GEN_5063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5065 = 9'h55 == r_count_12_io_out ? io_r_85_b : _GEN_5064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5066 = 9'h56 == r_count_12_io_out ? io_r_86_b : _GEN_5065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5067 = 9'h57 == r_count_12_io_out ? io_r_87_b : _GEN_5066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5068 = 9'h58 == r_count_12_io_out ? io_r_88_b : _GEN_5067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5069 = 9'h59 == r_count_12_io_out ? io_r_89_b : _GEN_5068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5070 = 9'h5a == r_count_12_io_out ? io_r_90_b : _GEN_5069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5071 = 9'h5b == r_count_12_io_out ? io_r_91_b : _GEN_5070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5072 = 9'h5c == r_count_12_io_out ? io_r_92_b : _GEN_5071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5073 = 9'h5d == r_count_12_io_out ? io_r_93_b : _GEN_5072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5074 = 9'h5e == r_count_12_io_out ? io_r_94_b : _GEN_5073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5075 = 9'h5f == r_count_12_io_out ? io_r_95_b : _GEN_5074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5076 = 9'h60 == r_count_12_io_out ? io_r_96_b : _GEN_5075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5077 = 9'h61 == r_count_12_io_out ? io_r_97_b : _GEN_5076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5078 = 9'h62 == r_count_12_io_out ? io_r_98_b : _GEN_5077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5079 = 9'h63 == r_count_12_io_out ? io_r_99_b : _GEN_5078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5080 = 9'h64 == r_count_12_io_out ? io_r_100_b : _GEN_5079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5081 = 9'h65 == r_count_12_io_out ? io_r_101_b : _GEN_5080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5082 = 9'h66 == r_count_12_io_out ? io_r_102_b : _GEN_5081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5083 = 9'h67 == r_count_12_io_out ? io_r_103_b : _GEN_5082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5084 = 9'h68 == r_count_12_io_out ? io_r_104_b : _GEN_5083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5085 = 9'h69 == r_count_12_io_out ? io_r_105_b : _GEN_5084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5086 = 9'h6a == r_count_12_io_out ? io_r_106_b : _GEN_5085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5087 = 9'h6b == r_count_12_io_out ? io_r_107_b : _GEN_5086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5088 = 9'h6c == r_count_12_io_out ? io_r_108_b : _GEN_5087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5089 = 9'h6d == r_count_12_io_out ? io_r_109_b : _GEN_5088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5090 = 9'h6e == r_count_12_io_out ? io_r_110_b : _GEN_5089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5091 = 9'h6f == r_count_12_io_out ? io_r_111_b : _GEN_5090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5092 = 9'h70 == r_count_12_io_out ? io_r_112_b : _GEN_5091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5093 = 9'h71 == r_count_12_io_out ? io_r_113_b : _GEN_5092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5094 = 9'h72 == r_count_12_io_out ? io_r_114_b : _GEN_5093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5095 = 9'h73 == r_count_12_io_out ? io_r_115_b : _GEN_5094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5096 = 9'h74 == r_count_12_io_out ? io_r_116_b : _GEN_5095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5097 = 9'h75 == r_count_12_io_out ? io_r_117_b : _GEN_5096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5098 = 9'h76 == r_count_12_io_out ? io_r_118_b : _GEN_5097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5099 = 9'h77 == r_count_12_io_out ? io_r_119_b : _GEN_5098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5100 = 9'h78 == r_count_12_io_out ? io_r_120_b : _GEN_5099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5101 = 9'h79 == r_count_12_io_out ? io_r_121_b : _GEN_5100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5102 = 9'h7a == r_count_12_io_out ? io_r_122_b : _GEN_5101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5103 = 9'h7b == r_count_12_io_out ? io_r_123_b : _GEN_5102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5104 = 9'h7c == r_count_12_io_out ? io_r_124_b : _GEN_5103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5105 = 9'h7d == r_count_12_io_out ? io_r_125_b : _GEN_5104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5106 = 9'h7e == r_count_12_io_out ? io_r_126_b : _GEN_5105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5107 = 9'h7f == r_count_12_io_out ? io_r_127_b : _GEN_5106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5108 = 9'h80 == r_count_12_io_out ? io_r_128_b : _GEN_5107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5109 = 9'h81 == r_count_12_io_out ? io_r_129_b : _GEN_5108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5110 = 9'h82 == r_count_12_io_out ? io_r_130_b : _GEN_5109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5111 = 9'h83 == r_count_12_io_out ? io_r_131_b : _GEN_5110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5112 = 9'h84 == r_count_12_io_out ? io_r_132_b : _GEN_5111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5113 = 9'h85 == r_count_12_io_out ? io_r_133_b : _GEN_5112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5114 = 9'h86 == r_count_12_io_out ? io_r_134_b : _GEN_5113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5115 = 9'h87 == r_count_12_io_out ? io_r_135_b : _GEN_5114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5116 = 9'h88 == r_count_12_io_out ? io_r_136_b : _GEN_5115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5117 = 9'h89 == r_count_12_io_out ? io_r_137_b : _GEN_5116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5118 = 9'h8a == r_count_12_io_out ? io_r_138_b : _GEN_5117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5119 = 9'h8b == r_count_12_io_out ? io_r_139_b : _GEN_5118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5120 = 9'h8c == r_count_12_io_out ? io_r_140_b : _GEN_5119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5121 = 9'h8d == r_count_12_io_out ? io_r_141_b : _GEN_5120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5122 = 9'h8e == r_count_12_io_out ? io_r_142_b : _GEN_5121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5123 = 9'h8f == r_count_12_io_out ? io_r_143_b : _GEN_5122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5124 = 9'h90 == r_count_12_io_out ? io_r_144_b : _GEN_5123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5125 = 9'h91 == r_count_12_io_out ? io_r_145_b : _GEN_5124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5126 = 9'h92 == r_count_12_io_out ? io_r_146_b : _GEN_5125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5127 = 9'h93 == r_count_12_io_out ? io_r_147_b : _GEN_5126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5128 = 9'h94 == r_count_12_io_out ? io_r_148_b : _GEN_5127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5129 = 9'h95 == r_count_12_io_out ? io_r_149_b : _GEN_5128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5130 = 9'h96 == r_count_12_io_out ? io_r_150_b : _GEN_5129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5131 = 9'h97 == r_count_12_io_out ? io_r_151_b : _GEN_5130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5132 = 9'h98 == r_count_12_io_out ? io_r_152_b : _GEN_5131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5133 = 9'h99 == r_count_12_io_out ? io_r_153_b : _GEN_5132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5134 = 9'h9a == r_count_12_io_out ? io_r_154_b : _GEN_5133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5135 = 9'h9b == r_count_12_io_out ? io_r_155_b : _GEN_5134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5136 = 9'h9c == r_count_12_io_out ? io_r_156_b : _GEN_5135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5137 = 9'h9d == r_count_12_io_out ? io_r_157_b : _GEN_5136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5138 = 9'h9e == r_count_12_io_out ? io_r_158_b : _GEN_5137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5139 = 9'h9f == r_count_12_io_out ? io_r_159_b : _GEN_5138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5140 = 9'ha0 == r_count_12_io_out ? io_r_160_b : _GEN_5139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5141 = 9'ha1 == r_count_12_io_out ? io_r_161_b : _GEN_5140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5142 = 9'ha2 == r_count_12_io_out ? io_r_162_b : _GEN_5141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5143 = 9'ha3 == r_count_12_io_out ? io_r_163_b : _GEN_5142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5144 = 9'ha4 == r_count_12_io_out ? io_r_164_b : _GEN_5143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5145 = 9'ha5 == r_count_12_io_out ? io_r_165_b : _GEN_5144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5146 = 9'ha6 == r_count_12_io_out ? io_r_166_b : _GEN_5145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5147 = 9'ha7 == r_count_12_io_out ? io_r_167_b : _GEN_5146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5148 = 9'ha8 == r_count_12_io_out ? io_r_168_b : _GEN_5147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5149 = 9'ha9 == r_count_12_io_out ? io_r_169_b : _GEN_5148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5150 = 9'haa == r_count_12_io_out ? io_r_170_b : _GEN_5149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5151 = 9'hab == r_count_12_io_out ? io_r_171_b : _GEN_5150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5152 = 9'hac == r_count_12_io_out ? io_r_172_b : _GEN_5151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5153 = 9'had == r_count_12_io_out ? io_r_173_b : _GEN_5152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5154 = 9'hae == r_count_12_io_out ? io_r_174_b : _GEN_5153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5155 = 9'haf == r_count_12_io_out ? io_r_175_b : _GEN_5154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5156 = 9'hb0 == r_count_12_io_out ? io_r_176_b : _GEN_5155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5157 = 9'hb1 == r_count_12_io_out ? io_r_177_b : _GEN_5156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5158 = 9'hb2 == r_count_12_io_out ? io_r_178_b : _GEN_5157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5159 = 9'hb3 == r_count_12_io_out ? io_r_179_b : _GEN_5158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5160 = 9'hb4 == r_count_12_io_out ? io_r_180_b : _GEN_5159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5161 = 9'hb5 == r_count_12_io_out ? io_r_181_b : _GEN_5160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5162 = 9'hb6 == r_count_12_io_out ? io_r_182_b : _GEN_5161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5163 = 9'hb7 == r_count_12_io_out ? io_r_183_b : _GEN_5162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5164 = 9'hb8 == r_count_12_io_out ? io_r_184_b : _GEN_5163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5165 = 9'hb9 == r_count_12_io_out ? io_r_185_b : _GEN_5164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5166 = 9'hba == r_count_12_io_out ? io_r_186_b : _GEN_5165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5167 = 9'hbb == r_count_12_io_out ? io_r_187_b : _GEN_5166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5168 = 9'hbc == r_count_12_io_out ? io_r_188_b : _GEN_5167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5169 = 9'hbd == r_count_12_io_out ? io_r_189_b : _GEN_5168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5170 = 9'hbe == r_count_12_io_out ? io_r_190_b : _GEN_5169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5171 = 9'hbf == r_count_12_io_out ? io_r_191_b : _GEN_5170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5172 = 9'hc0 == r_count_12_io_out ? io_r_192_b : _GEN_5171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5173 = 9'hc1 == r_count_12_io_out ? io_r_193_b : _GEN_5172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5174 = 9'hc2 == r_count_12_io_out ? io_r_194_b : _GEN_5173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5175 = 9'hc3 == r_count_12_io_out ? io_r_195_b : _GEN_5174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5176 = 9'hc4 == r_count_12_io_out ? io_r_196_b : _GEN_5175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5177 = 9'hc5 == r_count_12_io_out ? io_r_197_b : _GEN_5176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5178 = 9'hc6 == r_count_12_io_out ? io_r_198_b : _GEN_5177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5179 = 9'hc7 == r_count_12_io_out ? io_r_199_b : _GEN_5178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5180 = 9'hc8 == r_count_12_io_out ? io_r_200_b : _GEN_5179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5181 = 9'hc9 == r_count_12_io_out ? io_r_201_b : _GEN_5180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5182 = 9'hca == r_count_12_io_out ? io_r_202_b : _GEN_5181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5183 = 9'hcb == r_count_12_io_out ? io_r_203_b : _GEN_5182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5184 = 9'hcc == r_count_12_io_out ? io_r_204_b : _GEN_5183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5185 = 9'hcd == r_count_12_io_out ? io_r_205_b : _GEN_5184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5186 = 9'hce == r_count_12_io_out ? io_r_206_b : _GEN_5185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5187 = 9'hcf == r_count_12_io_out ? io_r_207_b : _GEN_5186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5188 = 9'hd0 == r_count_12_io_out ? io_r_208_b : _GEN_5187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5189 = 9'hd1 == r_count_12_io_out ? io_r_209_b : _GEN_5188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5190 = 9'hd2 == r_count_12_io_out ? io_r_210_b : _GEN_5189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5191 = 9'hd3 == r_count_12_io_out ? io_r_211_b : _GEN_5190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5192 = 9'hd4 == r_count_12_io_out ? io_r_212_b : _GEN_5191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5193 = 9'hd5 == r_count_12_io_out ? io_r_213_b : _GEN_5192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5194 = 9'hd6 == r_count_12_io_out ? io_r_214_b : _GEN_5193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5195 = 9'hd7 == r_count_12_io_out ? io_r_215_b : _GEN_5194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5196 = 9'hd8 == r_count_12_io_out ? io_r_216_b : _GEN_5195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5197 = 9'hd9 == r_count_12_io_out ? io_r_217_b : _GEN_5196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5198 = 9'hda == r_count_12_io_out ? io_r_218_b : _GEN_5197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5199 = 9'hdb == r_count_12_io_out ? io_r_219_b : _GEN_5198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5200 = 9'hdc == r_count_12_io_out ? io_r_220_b : _GEN_5199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5201 = 9'hdd == r_count_12_io_out ? io_r_221_b : _GEN_5200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5202 = 9'hde == r_count_12_io_out ? io_r_222_b : _GEN_5201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5203 = 9'hdf == r_count_12_io_out ? io_r_223_b : _GEN_5202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5204 = 9'he0 == r_count_12_io_out ? io_r_224_b : _GEN_5203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5205 = 9'he1 == r_count_12_io_out ? io_r_225_b : _GEN_5204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5206 = 9'he2 == r_count_12_io_out ? io_r_226_b : _GEN_5205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5207 = 9'he3 == r_count_12_io_out ? io_r_227_b : _GEN_5206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5208 = 9'he4 == r_count_12_io_out ? io_r_228_b : _GEN_5207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5209 = 9'he5 == r_count_12_io_out ? io_r_229_b : _GEN_5208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5210 = 9'he6 == r_count_12_io_out ? io_r_230_b : _GEN_5209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5211 = 9'he7 == r_count_12_io_out ? io_r_231_b : _GEN_5210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5212 = 9'he8 == r_count_12_io_out ? io_r_232_b : _GEN_5211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5213 = 9'he9 == r_count_12_io_out ? io_r_233_b : _GEN_5212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5214 = 9'hea == r_count_12_io_out ? io_r_234_b : _GEN_5213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5215 = 9'heb == r_count_12_io_out ? io_r_235_b : _GEN_5214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5216 = 9'hec == r_count_12_io_out ? io_r_236_b : _GEN_5215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5217 = 9'hed == r_count_12_io_out ? io_r_237_b : _GEN_5216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5218 = 9'hee == r_count_12_io_out ? io_r_238_b : _GEN_5217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5219 = 9'hef == r_count_12_io_out ? io_r_239_b : _GEN_5218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5220 = 9'hf0 == r_count_12_io_out ? io_r_240_b : _GEN_5219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5221 = 9'hf1 == r_count_12_io_out ? io_r_241_b : _GEN_5220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5222 = 9'hf2 == r_count_12_io_out ? io_r_242_b : _GEN_5221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5223 = 9'hf3 == r_count_12_io_out ? io_r_243_b : _GEN_5222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5224 = 9'hf4 == r_count_12_io_out ? io_r_244_b : _GEN_5223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5225 = 9'hf5 == r_count_12_io_out ? io_r_245_b : _GEN_5224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5226 = 9'hf6 == r_count_12_io_out ? io_r_246_b : _GEN_5225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5227 = 9'hf7 == r_count_12_io_out ? io_r_247_b : _GEN_5226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5228 = 9'hf8 == r_count_12_io_out ? io_r_248_b : _GEN_5227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5229 = 9'hf9 == r_count_12_io_out ? io_r_249_b : _GEN_5228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5230 = 9'hfa == r_count_12_io_out ? io_r_250_b : _GEN_5229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5231 = 9'hfb == r_count_12_io_out ? io_r_251_b : _GEN_5230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5232 = 9'hfc == r_count_12_io_out ? io_r_252_b : _GEN_5231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5233 = 9'hfd == r_count_12_io_out ? io_r_253_b : _GEN_5232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5234 = 9'hfe == r_count_12_io_out ? io_r_254_b : _GEN_5233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5235 = 9'hff == r_count_12_io_out ? io_r_255_b : _GEN_5234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5236 = 9'h100 == r_count_12_io_out ? io_r_256_b : _GEN_5235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5237 = 9'h101 == r_count_12_io_out ? io_r_257_b : _GEN_5236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5238 = 9'h102 == r_count_12_io_out ? io_r_258_b : _GEN_5237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5239 = 9'h103 == r_count_12_io_out ? io_r_259_b : _GEN_5238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5240 = 9'h104 == r_count_12_io_out ? io_r_260_b : _GEN_5239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5241 = 9'h105 == r_count_12_io_out ? io_r_261_b : _GEN_5240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5242 = 9'h106 == r_count_12_io_out ? io_r_262_b : _GEN_5241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5243 = 9'h107 == r_count_12_io_out ? io_r_263_b : _GEN_5242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5244 = 9'h108 == r_count_12_io_out ? io_r_264_b : _GEN_5243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5245 = 9'h109 == r_count_12_io_out ? io_r_265_b : _GEN_5244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5246 = 9'h10a == r_count_12_io_out ? io_r_266_b : _GEN_5245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5247 = 9'h10b == r_count_12_io_out ? io_r_267_b : _GEN_5246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5248 = 9'h10c == r_count_12_io_out ? io_r_268_b : _GEN_5247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5249 = 9'h10d == r_count_12_io_out ? io_r_269_b : _GEN_5248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5250 = 9'h10e == r_count_12_io_out ? io_r_270_b : _GEN_5249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5251 = 9'h10f == r_count_12_io_out ? io_r_271_b : _GEN_5250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5252 = 9'h110 == r_count_12_io_out ? io_r_272_b : _GEN_5251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5253 = 9'h111 == r_count_12_io_out ? io_r_273_b : _GEN_5252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5254 = 9'h112 == r_count_12_io_out ? io_r_274_b : _GEN_5253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5255 = 9'h113 == r_count_12_io_out ? io_r_275_b : _GEN_5254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5256 = 9'h114 == r_count_12_io_out ? io_r_276_b : _GEN_5255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5257 = 9'h115 == r_count_12_io_out ? io_r_277_b : _GEN_5256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5258 = 9'h116 == r_count_12_io_out ? io_r_278_b : _GEN_5257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5259 = 9'h117 == r_count_12_io_out ? io_r_279_b : _GEN_5258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5260 = 9'h118 == r_count_12_io_out ? io_r_280_b : _GEN_5259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5261 = 9'h119 == r_count_12_io_out ? io_r_281_b : _GEN_5260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5262 = 9'h11a == r_count_12_io_out ? io_r_282_b : _GEN_5261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5263 = 9'h11b == r_count_12_io_out ? io_r_283_b : _GEN_5262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5264 = 9'h11c == r_count_12_io_out ? io_r_284_b : _GEN_5263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5265 = 9'h11d == r_count_12_io_out ? io_r_285_b : _GEN_5264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5266 = 9'h11e == r_count_12_io_out ? io_r_286_b : _GEN_5265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5267 = 9'h11f == r_count_12_io_out ? io_r_287_b : _GEN_5266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5268 = 9'h120 == r_count_12_io_out ? io_r_288_b : _GEN_5267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5269 = 9'h121 == r_count_12_io_out ? io_r_289_b : _GEN_5268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5270 = 9'h122 == r_count_12_io_out ? io_r_290_b : _GEN_5269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5271 = 9'h123 == r_count_12_io_out ? io_r_291_b : _GEN_5270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5272 = 9'h124 == r_count_12_io_out ? io_r_292_b : _GEN_5271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5273 = 9'h125 == r_count_12_io_out ? io_r_293_b : _GEN_5272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5274 = 9'h126 == r_count_12_io_out ? io_r_294_b : _GEN_5273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5275 = 9'h127 == r_count_12_io_out ? io_r_295_b : _GEN_5274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5276 = 9'h128 == r_count_12_io_out ? io_r_296_b : _GEN_5275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5277 = 9'h129 == r_count_12_io_out ? io_r_297_b : _GEN_5276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5278 = 9'h12a == r_count_12_io_out ? io_r_298_b : _GEN_5277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5279 = 9'h12b == r_count_12_io_out ? io_r_299_b : _GEN_5278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5280 = 9'h12c == r_count_12_io_out ? io_r_300_b : _GEN_5279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5281 = 9'h12d == r_count_12_io_out ? io_r_301_b : _GEN_5280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5282 = 9'h12e == r_count_12_io_out ? io_r_302_b : _GEN_5281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5283 = 9'h12f == r_count_12_io_out ? io_r_303_b : _GEN_5282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5284 = 9'h130 == r_count_12_io_out ? io_r_304_b : _GEN_5283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5285 = 9'h131 == r_count_12_io_out ? io_r_305_b : _GEN_5284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5286 = 9'h132 == r_count_12_io_out ? io_r_306_b : _GEN_5285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5287 = 9'h133 == r_count_12_io_out ? io_r_307_b : _GEN_5286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5288 = 9'h134 == r_count_12_io_out ? io_r_308_b : _GEN_5287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5289 = 9'h135 == r_count_12_io_out ? io_r_309_b : _GEN_5288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5290 = 9'h136 == r_count_12_io_out ? io_r_310_b : _GEN_5289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5291 = 9'h137 == r_count_12_io_out ? io_r_311_b : _GEN_5290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5292 = 9'h138 == r_count_12_io_out ? io_r_312_b : _GEN_5291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5293 = 9'h139 == r_count_12_io_out ? io_r_313_b : _GEN_5292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5294 = 9'h13a == r_count_12_io_out ? io_r_314_b : _GEN_5293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5295 = 9'h13b == r_count_12_io_out ? io_r_315_b : _GEN_5294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5296 = 9'h13c == r_count_12_io_out ? io_r_316_b : _GEN_5295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5297 = 9'h13d == r_count_12_io_out ? io_r_317_b : _GEN_5296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5298 = 9'h13e == r_count_12_io_out ? io_r_318_b : _GEN_5297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5299 = 9'h13f == r_count_12_io_out ? io_r_319_b : _GEN_5298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5300 = 9'h140 == r_count_12_io_out ? io_r_320_b : _GEN_5299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5301 = 9'h141 == r_count_12_io_out ? io_r_321_b : _GEN_5300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5302 = 9'h142 == r_count_12_io_out ? io_r_322_b : _GEN_5301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5303 = 9'h143 == r_count_12_io_out ? io_r_323_b : _GEN_5302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5304 = 9'h144 == r_count_12_io_out ? io_r_324_b : _GEN_5303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5305 = 9'h145 == r_count_12_io_out ? io_r_325_b : _GEN_5304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5306 = 9'h146 == r_count_12_io_out ? io_r_326_b : _GEN_5305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5307 = 9'h147 == r_count_12_io_out ? io_r_327_b : _GEN_5306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5308 = 9'h148 == r_count_12_io_out ? io_r_328_b : _GEN_5307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5309 = 9'h149 == r_count_12_io_out ? io_r_329_b : _GEN_5308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5310 = 9'h14a == r_count_12_io_out ? io_r_330_b : _GEN_5309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5311 = 9'h14b == r_count_12_io_out ? io_r_331_b : _GEN_5310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5312 = 9'h14c == r_count_12_io_out ? io_r_332_b : _GEN_5311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5313 = 9'h14d == r_count_12_io_out ? io_r_333_b : _GEN_5312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5314 = 9'h14e == r_count_12_io_out ? io_r_334_b : _GEN_5313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5315 = 9'h14f == r_count_12_io_out ? io_r_335_b : _GEN_5314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5316 = 9'h150 == r_count_12_io_out ? io_r_336_b : _GEN_5315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5317 = 9'h151 == r_count_12_io_out ? io_r_337_b : _GEN_5316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5318 = 9'h152 == r_count_12_io_out ? io_r_338_b : _GEN_5317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5319 = 9'h153 == r_count_12_io_out ? io_r_339_b : _GEN_5318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5320 = 9'h154 == r_count_12_io_out ? io_r_340_b : _GEN_5319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5321 = 9'h155 == r_count_12_io_out ? io_r_341_b : _GEN_5320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5322 = 9'h156 == r_count_12_io_out ? io_r_342_b : _GEN_5321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5323 = 9'h157 == r_count_12_io_out ? io_r_343_b : _GEN_5322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5324 = 9'h158 == r_count_12_io_out ? io_r_344_b : _GEN_5323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5325 = 9'h159 == r_count_12_io_out ? io_r_345_b : _GEN_5324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5326 = 9'h15a == r_count_12_io_out ? io_r_346_b : _GEN_5325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5327 = 9'h15b == r_count_12_io_out ? io_r_347_b : _GEN_5326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5328 = 9'h15c == r_count_12_io_out ? io_r_348_b : _GEN_5327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5329 = 9'h15d == r_count_12_io_out ? io_r_349_b : _GEN_5328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5330 = 9'h15e == r_count_12_io_out ? io_r_350_b : _GEN_5329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5331 = 9'h15f == r_count_12_io_out ? io_r_351_b : _GEN_5330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5332 = 9'h160 == r_count_12_io_out ? io_r_352_b : _GEN_5331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5333 = 9'h161 == r_count_12_io_out ? io_r_353_b : _GEN_5332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5334 = 9'h162 == r_count_12_io_out ? io_r_354_b : _GEN_5333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5335 = 9'h163 == r_count_12_io_out ? io_r_355_b : _GEN_5334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5336 = 9'h164 == r_count_12_io_out ? io_r_356_b : _GEN_5335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5337 = 9'h165 == r_count_12_io_out ? io_r_357_b : _GEN_5336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5338 = 9'h166 == r_count_12_io_out ? io_r_358_b : _GEN_5337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5339 = 9'h167 == r_count_12_io_out ? io_r_359_b : _GEN_5338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5340 = 9'h168 == r_count_12_io_out ? io_r_360_b : _GEN_5339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5341 = 9'h169 == r_count_12_io_out ? io_r_361_b : _GEN_5340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5342 = 9'h16a == r_count_12_io_out ? io_r_362_b : _GEN_5341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5343 = 9'h16b == r_count_12_io_out ? io_r_363_b : _GEN_5342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5344 = 9'h16c == r_count_12_io_out ? io_r_364_b : _GEN_5343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5345 = 9'h16d == r_count_12_io_out ? io_r_365_b : _GEN_5344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5346 = 9'h16e == r_count_12_io_out ? io_r_366_b : _GEN_5345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5347 = 9'h16f == r_count_12_io_out ? io_r_367_b : _GEN_5346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5348 = 9'h170 == r_count_12_io_out ? io_r_368_b : _GEN_5347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5349 = 9'h171 == r_count_12_io_out ? io_r_369_b : _GEN_5348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5350 = 9'h172 == r_count_12_io_out ? io_r_370_b : _GEN_5349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5351 = 9'h173 == r_count_12_io_out ? io_r_371_b : _GEN_5350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5352 = 9'h174 == r_count_12_io_out ? io_r_372_b : _GEN_5351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5353 = 9'h175 == r_count_12_io_out ? io_r_373_b : _GEN_5352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5354 = 9'h176 == r_count_12_io_out ? io_r_374_b : _GEN_5353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5355 = 9'h177 == r_count_12_io_out ? io_r_375_b : _GEN_5354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5356 = 9'h178 == r_count_12_io_out ? io_r_376_b : _GEN_5355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5357 = 9'h179 == r_count_12_io_out ? io_r_377_b : _GEN_5356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5358 = 9'h17a == r_count_12_io_out ? io_r_378_b : _GEN_5357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5359 = 9'h17b == r_count_12_io_out ? io_r_379_b : _GEN_5358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5360 = 9'h17c == r_count_12_io_out ? io_r_380_b : _GEN_5359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5361 = 9'h17d == r_count_12_io_out ? io_r_381_b : _GEN_5360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5362 = 9'h17e == r_count_12_io_out ? io_r_382_b : _GEN_5361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5363 = 9'h17f == r_count_12_io_out ? io_r_383_b : _GEN_5362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5364 = 9'h180 == r_count_12_io_out ? io_r_384_b : _GEN_5363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5365 = 9'h181 == r_count_12_io_out ? io_r_385_b : _GEN_5364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5366 = 9'h182 == r_count_12_io_out ? io_r_386_b : _GEN_5365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5367 = 9'h183 == r_count_12_io_out ? io_r_387_b : _GEN_5366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5368 = 9'h184 == r_count_12_io_out ? io_r_388_b : _GEN_5367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5369 = 9'h185 == r_count_12_io_out ? io_r_389_b : _GEN_5368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5370 = 9'h186 == r_count_12_io_out ? io_r_390_b : _GEN_5369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5371 = 9'h187 == r_count_12_io_out ? io_r_391_b : _GEN_5370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5372 = 9'h188 == r_count_12_io_out ? io_r_392_b : _GEN_5371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5373 = 9'h189 == r_count_12_io_out ? io_r_393_b : _GEN_5372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5374 = 9'h18a == r_count_12_io_out ? io_r_394_b : _GEN_5373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5375 = 9'h18b == r_count_12_io_out ? io_r_395_b : _GEN_5374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5376 = 9'h18c == r_count_12_io_out ? io_r_396_b : _GEN_5375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5377 = 9'h18d == r_count_12_io_out ? io_r_397_b : _GEN_5376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5378 = 9'h18e == r_count_12_io_out ? io_r_398_b : _GEN_5377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5381 = 9'h1 == r_count_13_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5382 = 9'h2 == r_count_13_io_out ? io_r_2_b : _GEN_5381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5383 = 9'h3 == r_count_13_io_out ? io_r_3_b : _GEN_5382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5384 = 9'h4 == r_count_13_io_out ? io_r_4_b : _GEN_5383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5385 = 9'h5 == r_count_13_io_out ? io_r_5_b : _GEN_5384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5386 = 9'h6 == r_count_13_io_out ? io_r_6_b : _GEN_5385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5387 = 9'h7 == r_count_13_io_out ? io_r_7_b : _GEN_5386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5388 = 9'h8 == r_count_13_io_out ? io_r_8_b : _GEN_5387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5389 = 9'h9 == r_count_13_io_out ? io_r_9_b : _GEN_5388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5390 = 9'ha == r_count_13_io_out ? io_r_10_b : _GEN_5389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5391 = 9'hb == r_count_13_io_out ? io_r_11_b : _GEN_5390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5392 = 9'hc == r_count_13_io_out ? io_r_12_b : _GEN_5391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5393 = 9'hd == r_count_13_io_out ? io_r_13_b : _GEN_5392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5394 = 9'he == r_count_13_io_out ? io_r_14_b : _GEN_5393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5395 = 9'hf == r_count_13_io_out ? io_r_15_b : _GEN_5394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5396 = 9'h10 == r_count_13_io_out ? io_r_16_b : _GEN_5395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5397 = 9'h11 == r_count_13_io_out ? io_r_17_b : _GEN_5396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5398 = 9'h12 == r_count_13_io_out ? io_r_18_b : _GEN_5397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5399 = 9'h13 == r_count_13_io_out ? io_r_19_b : _GEN_5398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5400 = 9'h14 == r_count_13_io_out ? io_r_20_b : _GEN_5399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5401 = 9'h15 == r_count_13_io_out ? io_r_21_b : _GEN_5400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5402 = 9'h16 == r_count_13_io_out ? io_r_22_b : _GEN_5401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5403 = 9'h17 == r_count_13_io_out ? io_r_23_b : _GEN_5402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5404 = 9'h18 == r_count_13_io_out ? io_r_24_b : _GEN_5403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5405 = 9'h19 == r_count_13_io_out ? io_r_25_b : _GEN_5404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5406 = 9'h1a == r_count_13_io_out ? io_r_26_b : _GEN_5405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5407 = 9'h1b == r_count_13_io_out ? io_r_27_b : _GEN_5406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5408 = 9'h1c == r_count_13_io_out ? io_r_28_b : _GEN_5407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5409 = 9'h1d == r_count_13_io_out ? io_r_29_b : _GEN_5408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5410 = 9'h1e == r_count_13_io_out ? io_r_30_b : _GEN_5409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5411 = 9'h1f == r_count_13_io_out ? io_r_31_b : _GEN_5410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5412 = 9'h20 == r_count_13_io_out ? io_r_32_b : _GEN_5411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5413 = 9'h21 == r_count_13_io_out ? io_r_33_b : _GEN_5412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5414 = 9'h22 == r_count_13_io_out ? io_r_34_b : _GEN_5413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5415 = 9'h23 == r_count_13_io_out ? io_r_35_b : _GEN_5414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5416 = 9'h24 == r_count_13_io_out ? io_r_36_b : _GEN_5415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5417 = 9'h25 == r_count_13_io_out ? io_r_37_b : _GEN_5416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5418 = 9'h26 == r_count_13_io_out ? io_r_38_b : _GEN_5417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5419 = 9'h27 == r_count_13_io_out ? io_r_39_b : _GEN_5418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5420 = 9'h28 == r_count_13_io_out ? io_r_40_b : _GEN_5419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5421 = 9'h29 == r_count_13_io_out ? io_r_41_b : _GEN_5420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5422 = 9'h2a == r_count_13_io_out ? io_r_42_b : _GEN_5421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5423 = 9'h2b == r_count_13_io_out ? io_r_43_b : _GEN_5422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5424 = 9'h2c == r_count_13_io_out ? io_r_44_b : _GEN_5423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5425 = 9'h2d == r_count_13_io_out ? io_r_45_b : _GEN_5424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5426 = 9'h2e == r_count_13_io_out ? io_r_46_b : _GEN_5425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5427 = 9'h2f == r_count_13_io_out ? io_r_47_b : _GEN_5426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5428 = 9'h30 == r_count_13_io_out ? io_r_48_b : _GEN_5427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5429 = 9'h31 == r_count_13_io_out ? io_r_49_b : _GEN_5428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5430 = 9'h32 == r_count_13_io_out ? io_r_50_b : _GEN_5429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5431 = 9'h33 == r_count_13_io_out ? io_r_51_b : _GEN_5430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5432 = 9'h34 == r_count_13_io_out ? io_r_52_b : _GEN_5431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5433 = 9'h35 == r_count_13_io_out ? io_r_53_b : _GEN_5432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5434 = 9'h36 == r_count_13_io_out ? io_r_54_b : _GEN_5433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5435 = 9'h37 == r_count_13_io_out ? io_r_55_b : _GEN_5434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5436 = 9'h38 == r_count_13_io_out ? io_r_56_b : _GEN_5435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5437 = 9'h39 == r_count_13_io_out ? io_r_57_b : _GEN_5436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5438 = 9'h3a == r_count_13_io_out ? io_r_58_b : _GEN_5437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5439 = 9'h3b == r_count_13_io_out ? io_r_59_b : _GEN_5438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5440 = 9'h3c == r_count_13_io_out ? io_r_60_b : _GEN_5439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5441 = 9'h3d == r_count_13_io_out ? io_r_61_b : _GEN_5440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5442 = 9'h3e == r_count_13_io_out ? io_r_62_b : _GEN_5441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5443 = 9'h3f == r_count_13_io_out ? io_r_63_b : _GEN_5442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5444 = 9'h40 == r_count_13_io_out ? io_r_64_b : _GEN_5443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5445 = 9'h41 == r_count_13_io_out ? io_r_65_b : _GEN_5444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5446 = 9'h42 == r_count_13_io_out ? io_r_66_b : _GEN_5445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5447 = 9'h43 == r_count_13_io_out ? io_r_67_b : _GEN_5446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5448 = 9'h44 == r_count_13_io_out ? io_r_68_b : _GEN_5447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5449 = 9'h45 == r_count_13_io_out ? io_r_69_b : _GEN_5448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5450 = 9'h46 == r_count_13_io_out ? io_r_70_b : _GEN_5449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5451 = 9'h47 == r_count_13_io_out ? io_r_71_b : _GEN_5450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5452 = 9'h48 == r_count_13_io_out ? io_r_72_b : _GEN_5451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5453 = 9'h49 == r_count_13_io_out ? io_r_73_b : _GEN_5452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5454 = 9'h4a == r_count_13_io_out ? io_r_74_b : _GEN_5453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5455 = 9'h4b == r_count_13_io_out ? io_r_75_b : _GEN_5454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5456 = 9'h4c == r_count_13_io_out ? io_r_76_b : _GEN_5455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5457 = 9'h4d == r_count_13_io_out ? io_r_77_b : _GEN_5456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5458 = 9'h4e == r_count_13_io_out ? io_r_78_b : _GEN_5457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5459 = 9'h4f == r_count_13_io_out ? io_r_79_b : _GEN_5458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5460 = 9'h50 == r_count_13_io_out ? io_r_80_b : _GEN_5459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5461 = 9'h51 == r_count_13_io_out ? io_r_81_b : _GEN_5460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5462 = 9'h52 == r_count_13_io_out ? io_r_82_b : _GEN_5461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5463 = 9'h53 == r_count_13_io_out ? io_r_83_b : _GEN_5462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5464 = 9'h54 == r_count_13_io_out ? io_r_84_b : _GEN_5463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5465 = 9'h55 == r_count_13_io_out ? io_r_85_b : _GEN_5464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5466 = 9'h56 == r_count_13_io_out ? io_r_86_b : _GEN_5465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5467 = 9'h57 == r_count_13_io_out ? io_r_87_b : _GEN_5466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5468 = 9'h58 == r_count_13_io_out ? io_r_88_b : _GEN_5467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5469 = 9'h59 == r_count_13_io_out ? io_r_89_b : _GEN_5468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5470 = 9'h5a == r_count_13_io_out ? io_r_90_b : _GEN_5469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5471 = 9'h5b == r_count_13_io_out ? io_r_91_b : _GEN_5470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5472 = 9'h5c == r_count_13_io_out ? io_r_92_b : _GEN_5471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5473 = 9'h5d == r_count_13_io_out ? io_r_93_b : _GEN_5472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5474 = 9'h5e == r_count_13_io_out ? io_r_94_b : _GEN_5473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5475 = 9'h5f == r_count_13_io_out ? io_r_95_b : _GEN_5474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5476 = 9'h60 == r_count_13_io_out ? io_r_96_b : _GEN_5475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5477 = 9'h61 == r_count_13_io_out ? io_r_97_b : _GEN_5476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5478 = 9'h62 == r_count_13_io_out ? io_r_98_b : _GEN_5477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5479 = 9'h63 == r_count_13_io_out ? io_r_99_b : _GEN_5478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5480 = 9'h64 == r_count_13_io_out ? io_r_100_b : _GEN_5479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5481 = 9'h65 == r_count_13_io_out ? io_r_101_b : _GEN_5480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5482 = 9'h66 == r_count_13_io_out ? io_r_102_b : _GEN_5481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5483 = 9'h67 == r_count_13_io_out ? io_r_103_b : _GEN_5482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5484 = 9'h68 == r_count_13_io_out ? io_r_104_b : _GEN_5483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5485 = 9'h69 == r_count_13_io_out ? io_r_105_b : _GEN_5484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5486 = 9'h6a == r_count_13_io_out ? io_r_106_b : _GEN_5485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5487 = 9'h6b == r_count_13_io_out ? io_r_107_b : _GEN_5486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5488 = 9'h6c == r_count_13_io_out ? io_r_108_b : _GEN_5487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5489 = 9'h6d == r_count_13_io_out ? io_r_109_b : _GEN_5488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5490 = 9'h6e == r_count_13_io_out ? io_r_110_b : _GEN_5489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5491 = 9'h6f == r_count_13_io_out ? io_r_111_b : _GEN_5490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5492 = 9'h70 == r_count_13_io_out ? io_r_112_b : _GEN_5491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5493 = 9'h71 == r_count_13_io_out ? io_r_113_b : _GEN_5492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5494 = 9'h72 == r_count_13_io_out ? io_r_114_b : _GEN_5493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5495 = 9'h73 == r_count_13_io_out ? io_r_115_b : _GEN_5494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5496 = 9'h74 == r_count_13_io_out ? io_r_116_b : _GEN_5495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5497 = 9'h75 == r_count_13_io_out ? io_r_117_b : _GEN_5496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5498 = 9'h76 == r_count_13_io_out ? io_r_118_b : _GEN_5497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5499 = 9'h77 == r_count_13_io_out ? io_r_119_b : _GEN_5498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5500 = 9'h78 == r_count_13_io_out ? io_r_120_b : _GEN_5499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5501 = 9'h79 == r_count_13_io_out ? io_r_121_b : _GEN_5500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5502 = 9'h7a == r_count_13_io_out ? io_r_122_b : _GEN_5501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5503 = 9'h7b == r_count_13_io_out ? io_r_123_b : _GEN_5502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5504 = 9'h7c == r_count_13_io_out ? io_r_124_b : _GEN_5503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5505 = 9'h7d == r_count_13_io_out ? io_r_125_b : _GEN_5504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5506 = 9'h7e == r_count_13_io_out ? io_r_126_b : _GEN_5505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5507 = 9'h7f == r_count_13_io_out ? io_r_127_b : _GEN_5506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5508 = 9'h80 == r_count_13_io_out ? io_r_128_b : _GEN_5507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5509 = 9'h81 == r_count_13_io_out ? io_r_129_b : _GEN_5508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5510 = 9'h82 == r_count_13_io_out ? io_r_130_b : _GEN_5509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5511 = 9'h83 == r_count_13_io_out ? io_r_131_b : _GEN_5510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5512 = 9'h84 == r_count_13_io_out ? io_r_132_b : _GEN_5511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5513 = 9'h85 == r_count_13_io_out ? io_r_133_b : _GEN_5512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5514 = 9'h86 == r_count_13_io_out ? io_r_134_b : _GEN_5513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5515 = 9'h87 == r_count_13_io_out ? io_r_135_b : _GEN_5514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5516 = 9'h88 == r_count_13_io_out ? io_r_136_b : _GEN_5515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5517 = 9'h89 == r_count_13_io_out ? io_r_137_b : _GEN_5516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5518 = 9'h8a == r_count_13_io_out ? io_r_138_b : _GEN_5517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5519 = 9'h8b == r_count_13_io_out ? io_r_139_b : _GEN_5518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5520 = 9'h8c == r_count_13_io_out ? io_r_140_b : _GEN_5519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5521 = 9'h8d == r_count_13_io_out ? io_r_141_b : _GEN_5520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5522 = 9'h8e == r_count_13_io_out ? io_r_142_b : _GEN_5521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5523 = 9'h8f == r_count_13_io_out ? io_r_143_b : _GEN_5522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5524 = 9'h90 == r_count_13_io_out ? io_r_144_b : _GEN_5523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5525 = 9'h91 == r_count_13_io_out ? io_r_145_b : _GEN_5524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5526 = 9'h92 == r_count_13_io_out ? io_r_146_b : _GEN_5525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5527 = 9'h93 == r_count_13_io_out ? io_r_147_b : _GEN_5526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5528 = 9'h94 == r_count_13_io_out ? io_r_148_b : _GEN_5527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5529 = 9'h95 == r_count_13_io_out ? io_r_149_b : _GEN_5528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5530 = 9'h96 == r_count_13_io_out ? io_r_150_b : _GEN_5529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5531 = 9'h97 == r_count_13_io_out ? io_r_151_b : _GEN_5530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5532 = 9'h98 == r_count_13_io_out ? io_r_152_b : _GEN_5531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5533 = 9'h99 == r_count_13_io_out ? io_r_153_b : _GEN_5532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5534 = 9'h9a == r_count_13_io_out ? io_r_154_b : _GEN_5533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5535 = 9'h9b == r_count_13_io_out ? io_r_155_b : _GEN_5534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5536 = 9'h9c == r_count_13_io_out ? io_r_156_b : _GEN_5535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5537 = 9'h9d == r_count_13_io_out ? io_r_157_b : _GEN_5536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5538 = 9'h9e == r_count_13_io_out ? io_r_158_b : _GEN_5537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5539 = 9'h9f == r_count_13_io_out ? io_r_159_b : _GEN_5538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5540 = 9'ha0 == r_count_13_io_out ? io_r_160_b : _GEN_5539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5541 = 9'ha1 == r_count_13_io_out ? io_r_161_b : _GEN_5540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5542 = 9'ha2 == r_count_13_io_out ? io_r_162_b : _GEN_5541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5543 = 9'ha3 == r_count_13_io_out ? io_r_163_b : _GEN_5542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5544 = 9'ha4 == r_count_13_io_out ? io_r_164_b : _GEN_5543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5545 = 9'ha5 == r_count_13_io_out ? io_r_165_b : _GEN_5544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5546 = 9'ha6 == r_count_13_io_out ? io_r_166_b : _GEN_5545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5547 = 9'ha7 == r_count_13_io_out ? io_r_167_b : _GEN_5546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5548 = 9'ha8 == r_count_13_io_out ? io_r_168_b : _GEN_5547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5549 = 9'ha9 == r_count_13_io_out ? io_r_169_b : _GEN_5548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5550 = 9'haa == r_count_13_io_out ? io_r_170_b : _GEN_5549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5551 = 9'hab == r_count_13_io_out ? io_r_171_b : _GEN_5550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5552 = 9'hac == r_count_13_io_out ? io_r_172_b : _GEN_5551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5553 = 9'had == r_count_13_io_out ? io_r_173_b : _GEN_5552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5554 = 9'hae == r_count_13_io_out ? io_r_174_b : _GEN_5553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5555 = 9'haf == r_count_13_io_out ? io_r_175_b : _GEN_5554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5556 = 9'hb0 == r_count_13_io_out ? io_r_176_b : _GEN_5555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5557 = 9'hb1 == r_count_13_io_out ? io_r_177_b : _GEN_5556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5558 = 9'hb2 == r_count_13_io_out ? io_r_178_b : _GEN_5557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5559 = 9'hb3 == r_count_13_io_out ? io_r_179_b : _GEN_5558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5560 = 9'hb4 == r_count_13_io_out ? io_r_180_b : _GEN_5559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5561 = 9'hb5 == r_count_13_io_out ? io_r_181_b : _GEN_5560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5562 = 9'hb6 == r_count_13_io_out ? io_r_182_b : _GEN_5561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5563 = 9'hb7 == r_count_13_io_out ? io_r_183_b : _GEN_5562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5564 = 9'hb8 == r_count_13_io_out ? io_r_184_b : _GEN_5563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5565 = 9'hb9 == r_count_13_io_out ? io_r_185_b : _GEN_5564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5566 = 9'hba == r_count_13_io_out ? io_r_186_b : _GEN_5565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5567 = 9'hbb == r_count_13_io_out ? io_r_187_b : _GEN_5566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5568 = 9'hbc == r_count_13_io_out ? io_r_188_b : _GEN_5567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5569 = 9'hbd == r_count_13_io_out ? io_r_189_b : _GEN_5568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5570 = 9'hbe == r_count_13_io_out ? io_r_190_b : _GEN_5569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5571 = 9'hbf == r_count_13_io_out ? io_r_191_b : _GEN_5570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5572 = 9'hc0 == r_count_13_io_out ? io_r_192_b : _GEN_5571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5573 = 9'hc1 == r_count_13_io_out ? io_r_193_b : _GEN_5572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5574 = 9'hc2 == r_count_13_io_out ? io_r_194_b : _GEN_5573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5575 = 9'hc3 == r_count_13_io_out ? io_r_195_b : _GEN_5574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5576 = 9'hc4 == r_count_13_io_out ? io_r_196_b : _GEN_5575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5577 = 9'hc5 == r_count_13_io_out ? io_r_197_b : _GEN_5576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5578 = 9'hc6 == r_count_13_io_out ? io_r_198_b : _GEN_5577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5579 = 9'hc7 == r_count_13_io_out ? io_r_199_b : _GEN_5578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5580 = 9'hc8 == r_count_13_io_out ? io_r_200_b : _GEN_5579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5581 = 9'hc9 == r_count_13_io_out ? io_r_201_b : _GEN_5580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5582 = 9'hca == r_count_13_io_out ? io_r_202_b : _GEN_5581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5583 = 9'hcb == r_count_13_io_out ? io_r_203_b : _GEN_5582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5584 = 9'hcc == r_count_13_io_out ? io_r_204_b : _GEN_5583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5585 = 9'hcd == r_count_13_io_out ? io_r_205_b : _GEN_5584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5586 = 9'hce == r_count_13_io_out ? io_r_206_b : _GEN_5585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5587 = 9'hcf == r_count_13_io_out ? io_r_207_b : _GEN_5586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5588 = 9'hd0 == r_count_13_io_out ? io_r_208_b : _GEN_5587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5589 = 9'hd1 == r_count_13_io_out ? io_r_209_b : _GEN_5588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5590 = 9'hd2 == r_count_13_io_out ? io_r_210_b : _GEN_5589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5591 = 9'hd3 == r_count_13_io_out ? io_r_211_b : _GEN_5590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5592 = 9'hd4 == r_count_13_io_out ? io_r_212_b : _GEN_5591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5593 = 9'hd5 == r_count_13_io_out ? io_r_213_b : _GEN_5592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5594 = 9'hd6 == r_count_13_io_out ? io_r_214_b : _GEN_5593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5595 = 9'hd7 == r_count_13_io_out ? io_r_215_b : _GEN_5594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5596 = 9'hd8 == r_count_13_io_out ? io_r_216_b : _GEN_5595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5597 = 9'hd9 == r_count_13_io_out ? io_r_217_b : _GEN_5596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5598 = 9'hda == r_count_13_io_out ? io_r_218_b : _GEN_5597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5599 = 9'hdb == r_count_13_io_out ? io_r_219_b : _GEN_5598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5600 = 9'hdc == r_count_13_io_out ? io_r_220_b : _GEN_5599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5601 = 9'hdd == r_count_13_io_out ? io_r_221_b : _GEN_5600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5602 = 9'hde == r_count_13_io_out ? io_r_222_b : _GEN_5601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5603 = 9'hdf == r_count_13_io_out ? io_r_223_b : _GEN_5602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5604 = 9'he0 == r_count_13_io_out ? io_r_224_b : _GEN_5603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5605 = 9'he1 == r_count_13_io_out ? io_r_225_b : _GEN_5604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5606 = 9'he2 == r_count_13_io_out ? io_r_226_b : _GEN_5605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5607 = 9'he3 == r_count_13_io_out ? io_r_227_b : _GEN_5606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5608 = 9'he4 == r_count_13_io_out ? io_r_228_b : _GEN_5607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5609 = 9'he5 == r_count_13_io_out ? io_r_229_b : _GEN_5608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5610 = 9'he6 == r_count_13_io_out ? io_r_230_b : _GEN_5609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5611 = 9'he7 == r_count_13_io_out ? io_r_231_b : _GEN_5610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5612 = 9'he8 == r_count_13_io_out ? io_r_232_b : _GEN_5611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5613 = 9'he9 == r_count_13_io_out ? io_r_233_b : _GEN_5612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5614 = 9'hea == r_count_13_io_out ? io_r_234_b : _GEN_5613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5615 = 9'heb == r_count_13_io_out ? io_r_235_b : _GEN_5614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5616 = 9'hec == r_count_13_io_out ? io_r_236_b : _GEN_5615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5617 = 9'hed == r_count_13_io_out ? io_r_237_b : _GEN_5616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5618 = 9'hee == r_count_13_io_out ? io_r_238_b : _GEN_5617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5619 = 9'hef == r_count_13_io_out ? io_r_239_b : _GEN_5618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5620 = 9'hf0 == r_count_13_io_out ? io_r_240_b : _GEN_5619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5621 = 9'hf1 == r_count_13_io_out ? io_r_241_b : _GEN_5620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5622 = 9'hf2 == r_count_13_io_out ? io_r_242_b : _GEN_5621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5623 = 9'hf3 == r_count_13_io_out ? io_r_243_b : _GEN_5622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5624 = 9'hf4 == r_count_13_io_out ? io_r_244_b : _GEN_5623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5625 = 9'hf5 == r_count_13_io_out ? io_r_245_b : _GEN_5624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5626 = 9'hf6 == r_count_13_io_out ? io_r_246_b : _GEN_5625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5627 = 9'hf7 == r_count_13_io_out ? io_r_247_b : _GEN_5626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5628 = 9'hf8 == r_count_13_io_out ? io_r_248_b : _GEN_5627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5629 = 9'hf9 == r_count_13_io_out ? io_r_249_b : _GEN_5628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5630 = 9'hfa == r_count_13_io_out ? io_r_250_b : _GEN_5629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5631 = 9'hfb == r_count_13_io_out ? io_r_251_b : _GEN_5630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5632 = 9'hfc == r_count_13_io_out ? io_r_252_b : _GEN_5631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5633 = 9'hfd == r_count_13_io_out ? io_r_253_b : _GEN_5632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5634 = 9'hfe == r_count_13_io_out ? io_r_254_b : _GEN_5633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5635 = 9'hff == r_count_13_io_out ? io_r_255_b : _GEN_5634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5636 = 9'h100 == r_count_13_io_out ? io_r_256_b : _GEN_5635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5637 = 9'h101 == r_count_13_io_out ? io_r_257_b : _GEN_5636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5638 = 9'h102 == r_count_13_io_out ? io_r_258_b : _GEN_5637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5639 = 9'h103 == r_count_13_io_out ? io_r_259_b : _GEN_5638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5640 = 9'h104 == r_count_13_io_out ? io_r_260_b : _GEN_5639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5641 = 9'h105 == r_count_13_io_out ? io_r_261_b : _GEN_5640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5642 = 9'h106 == r_count_13_io_out ? io_r_262_b : _GEN_5641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5643 = 9'h107 == r_count_13_io_out ? io_r_263_b : _GEN_5642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5644 = 9'h108 == r_count_13_io_out ? io_r_264_b : _GEN_5643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5645 = 9'h109 == r_count_13_io_out ? io_r_265_b : _GEN_5644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5646 = 9'h10a == r_count_13_io_out ? io_r_266_b : _GEN_5645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5647 = 9'h10b == r_count_13_io_out ? io_r_267_b : _GEN_5646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5648 = 9'h10c == r_count_13_io_out ? io_r_268_b : _GEN_5647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5649 = 9'h10d == r_count_13_io_out ? io_r_269_b : _GEN_5648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5650 = 9'h10e == r_count_13_io_out ? io_r_270_b : _GEN_5649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5651 = 9'h10f == r_count_13_io_out ? io_r_271_b : _GEN_5650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5652 = 9'h110 == r_count_13_io_out ? io_r_272_b : _GEN_5651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5653 = 9'h111 == r_count_13_io_out ? io_r_273_b : _GEN_5652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5654 = 9'h112 == r_count_13_io_out ? io_r_274_b : _GEN_5653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5655 = 9'h113 == r_count_13_io_out ? io_r_275_b : _GEN_5654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5656 = 9'h114 == r_count_13_io_out ? io_r_276_b : _GEN_5655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5657 = 9'h115 == r_count_13_io_out ? io_r_277_b : _GEN_5656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5658 = 9'h116 == r_count_13_io_out ? io_r_278_b : _GEN_5657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5659 = 9'h117 == r_count_13_io_out ? io_r_279_b : _GEN_5658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5660 = 9'h118 == r_count_13_io_out ? io_r_280_b : _GEN_5659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5661 = 9'h119 == r_count_13_io_out ? io_r_281_b : _GEN_5660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5662 = 9'h11a == r_count_13_io_out ? io_r_282_b : _GEN_5661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5663 = 9'h11b == r_count_13_io_out ? io_r_283_b : _GEN_5662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5664 = 9'h11c == r_count_13_io_out ? io_r_284_b : _GEN_5663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5665 = 9'h11d == r_count_13_io_out ? io_r_285_b : _GEN_5664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5666 = 9'h11e == r_count_13_io_out ? io_r_286_b : _GEN_5665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5667 = 9'h11f == r_count_13_io_out ? io_r_287_b : _GEN_5666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5668 = 9'h120 == r_count_13_io_out ? io_r_288_b : _GEN_5667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5669 = 9'h121 == r_count_13_io_out ? io_r_289_b : _GEN_5668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5670 = 9'h122 == r_count_13_io_out ? io_r_290_b : _GEN_5669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5671 = 9'h123 == r_count_13_io_out ? io_r_291_b : _GEN_5670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5672 = 9'h124 == r_count_13_io_out ? io_r_292_b : _GEN_5671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5673 = 9'h125 == r_count_13_io_out ? io_r_293_b : _GEN_5672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5674 = 9'h126 == r_count_13_io_out ? io_r_294_b : _GEN_5673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5675 = 9'h127 == r_count_13_io_out ? io_r_295_b : _GEN_5674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5676 = 9'h128 == r_count_13_io_out ? io_r_296_b : _GEN_5675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5677 = 9'h129 == r_count_13_io_out ? io_r_297_b : _GEN_5676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5678 = 9'h12a == r_count_13_io_out ? io_r_298_b : _GEN_5677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5679 = 9'h12b == r_count_13_io_out ? io_r_299_b : _GEN_5678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5680 = 9'h12c == r_count_13_io_out ? io_r_300_b : _GEN_5679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5681 = 9'h12d == r_count_13_io_out ? io_r_301_b : _GEN_5680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5682 = 9'h12e == r_count_13_io_out ? io_r_302_b : _GEN_5681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5683 = 9'h12f == r_count_13_io_out ? io_r_303_b : _GEN_5682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5684 = 9'h130 == r_count_13_io_out ? io_r_304_b : _GEN_5683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5685 = 9'h131 == r_count_13_io_out ? io_r_305_b : _GEN_5684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5686 = 9'h132 == r_count_13_io_out ? io_r_306_b : _GEN_5685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5687 = 9'h133 == r_count_13_io_out ? io_r_307_b : _GEN_5686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5688 = 9'h134 == r_count_13_io_out ? io_r_308_b : _GEN_5687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5689 = 9'h135 == r_count_13_io_out ? io_r_309_b : _GEN_5688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5690 = 9'h136 == r_count_13_io_out ? io_r_310_b : _GEN_5689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5691 = 9'h137 == r_count_13_io_out ? io_r_311_b : _GEN_5690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5692 = 9'h138 == r_count_13_io_out ? io_r_312_b : _GEN_5691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5693 = 9'h139 == r_count_13_io_out ? io_r_313_b : _GEN_5692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5694 = 9'h13a == r_count_13_io_out ? io_r_314_b : _GEN_5693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5695 = 9'h13b == r_count_13_io_out ? io_r_315_b : _GEN_5694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5696 = 9'h13c == r_count_13_io_out ? io_r_316_b : _GEN_5695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5697 = 9'h13d == r_count_13_io_out ? io_r_317_b : _GEN_5696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5698 = 9'h13e == r_count_13_io_out ? io_r_318_b : _GEN_5697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5699 = 9'h13f == r_count_13_io_out ? io_r_319_b : _GEN_5698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5700 = 9'h140 == r_count_13_io_out ? io_r_320_b : _GEN_5699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5701 = 9'h141 == r_count_13_io_out ? io_r_321_b : _GEN_5700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5702 = 9'h142 == r_count_13_io_out ? io_r_322_b : _GEN_5701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5703 = 9'h143 == r_count_13_io_out ? io_r_323_b : _GEN_5702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5704 = 9'h144 == r_count_13_io_out ? io_r_324_b : _GEN_5703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5705 = 9'h145 == r_count_13_io_out ? io_r_325_b : _GEN_5704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5706 = 9'h146 == r_count_13_io_out ? io_r_326_b : _GEN_5705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5707 = 9'h147 == r_count_13_io_out ? io_r_327_b : _GEN_5706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5708 = 9'h148 == r_count_13_io_out ? io_r_328_b : _GEN_5707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5709 = 9'h149 == r_count_13_io_out ? io_r_329_b : _GEN_5708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5710 = 9'h14a == r_count_13_io_out ? io_r_330_b : _GEN_5709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5711 = 9'h14b == r_count_13_io_out ? io_r_331_b : _GEN_5710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5712 = 9'h14c == r_count_13_io_out ? io_r_332_b : _GEN_5711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5713 = 9'h14d == r_count_13_io_out ? io_r_333_b : _GEN_5712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5714 = 9'h14e == r_count_13_io_out ? io_r_334_b : _GEN_5713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5715 = 9'h14f == r_count_13_io_out ? io_r_335_b : _GEN_5714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5716 = 9'h150 == r_count_13_io_out ? io_r_336_b : _GEN_5715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5717 = 9'h151 == r_count_13_io_out ? io_r_337_b : _GEN_5716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5718 = 9'h152 == r_count_13_io_out ? io_r_338_b : _GEN_5717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5719 = 9'h153 == r_count_13_io_out ? io_r_339_b : _GEN_5718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5720 = 9'h154 == r_count_13_io_out ? io_r_340_b : _GEN_5719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5721 = 9'h155 == r_count_13_io_out ? io_r_341_b : _GEN_5720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5722 = 9'h156 == r_count_13_io_out ? io_r_342_b : _GEN_5721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5723 = 9'h157 == r_count_13_io_out ? io_r_343_b : _GEN_5722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5724 = 9'h158 == r_count_13_io_out ? io_r_344_b : _GEN_5723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5725 = 9'h159 == r_count_13_io_out ? io_r_345_b : _GEN_5724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5726 = 9'h15a == r_count_13_io_out ? io_r_346_b : _GEN_5725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5727 = 9'h15b == r_count_13_io_out ? io_r_347_b : _GEN_5726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5728 = 9'h15c == r_count_13_io_out ? io_r_348_b : _GEN_5727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5729 = 9'h15d == r_count_13_io_out ? io_r_349_b : _GEN_5728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5730 = 9'h15e == r_count_13_io_out ? io_r_350_b : _GEN_5729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5731 = 9'h15f == r_count_13_io_out ? io_r_351_b : _GEN_5730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5732 = 9'h160 == r_count_13_io_out ? io_r_352_b : _GEN_5731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5733 = 9'h161 == r_count_13_io_out ? io_r_353_b : _GEN_5732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5734 = 9'h162 == r_count_13_io_out ? io_r_354_b : _GEN_5733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5735 = 9'h163 == r_count_13_io_out ? io_r_355_b : _GEN_5734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5736 = 9'h164 == r_count_13_io_out ? io_r_356_b : _GEN_5735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5737 = 9'h165 == r_count_13_io_out ? io_r_357_b : _GEN_5736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5738 = 9'h166 == r_count_13_io_out ? io_r_358_b : _GEN_5737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5739 = 9'h167 == r_count_13_io_out ? io_r_359_b : _GEN_5738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5740 = 9'h168 == r_count_13_io_out ? io_r_360_b : _GEN_5739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5741 = 9'h169 == r_count_13_io_out ? io_r_361_b : _GEN_5740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5742 = 9'h16a == r_count_13_io_out ? io_r_362_b : _GEN_5741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5743 = 9'h16b == r_count_13_io_out ? io_r_363_b : _GEN_5742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5744 = 9'h16c == r_count_13_io_out ? io_r_364_b : _GEN_5743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5745 = 9'h16d == r_count_13_io_out ? io_r_365_b : _GEN_5744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5746 = 9'h16e == r_count_13_io_out ? io_r_366_b : _GEN_5745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5747 = 9'h16f == r_count_13_io_out ? io_r_367_b : _GEN_5746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5748 = 9'h170 == r_count_13_io_out ? io_r_368_b : _GEN_5747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5749 = 9'h171 == r_count_13_io_out ? io_r_369_b : _GEN_5748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5750 = 9'h172 == r_count_13_io_out ? io_r_370_b : _GEN_5749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5751 = 9'h173 == r_count_13_io_out ? io_r_371_b : _GEN_5750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5752 = 9'h174 == r_count_13_io_out ? io_r_372_b : _GEN_5751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5753 = 9'h175 == r_count_13_io_out ? io_r_373_b : _GEN_5752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5754 = 9'h176 == r_count_13_io_out ? io_r_374_b : _GEN_5753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5755 = 9'h177 == r_count_13_io_out ? io_r_375_b : _GEN_5754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5756 = 9'h178 == r_count_13_io_out ? io_r_376_b : _GEN_5755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5757 = 9'h179 == r_count_13_io_out ? io_r_377_b : _GEN_5756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5758 = 9'h17a == r_count_13_io_out ? io_r_378_b : _GEN_5757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5759 = 9'h17b == r_count_13_io_out ? io_r_379_b : _GEN_5758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5760 = 9'h17c == r_count_13_io_out ? io_r_380_b : _GEN_5759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5761 = 9'h17d == r_count_13_io_out ? io_r_381_b : _GEN_5760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5762 = 9'h17e == r_count_13_io_out ? io_r_382_b : _GEN_5761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5763 = 9'h17f == r_count_13_io_out ? io_r_383_b : _GEN_5762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5764 = 9'h180 == r_count_13_io_out ? io_r_384_b : _GEN_5763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5765 = 9'h181 == r_count_13_io_out ? io_r_385_b : _GEN_5764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5766 = 9'h182 == r_count_13_io_out ? io_r_386_b : _GEN_5765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5767 = 9'h183 == r_count_13_io_out ? io_r_387_b : _GEN_5766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5768 = 9'h184 == r_count_13_io_out ? io_r_388_b : _GEN_5767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5769 = 9'h185 == r_count_13_io_out ? io_r_389_b : _GEN_5768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5770 = 9'h186 == r_count_13_io_out ? io_r_390_b : _GEN_5769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5771 = 9'h187 == r_count_13_io_out ? io_r_391_b : _GEN_5770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5772 = 9'h188 == r_count_13_io_out ? io_r_392_b : _GEN_5771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5773 = 9'h189 == r_count_13_io_out ? io_r_393_b : _GEN_5772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5774 = 9'h18a == r_count_13_io_out ? io_r_394_b : _GEN_5773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5775 = 9'h18b == r_count_13_io_out ? io_r_395_b : _GEN_5774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5776 = 9'h18c == r_count_13_io_out ? io_r_396_b : _GEN_5775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5777 = 9'h18d == r_count_13_io_out ? io_r_397_b : _GEN_5776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5778 = 9'h18e == r_count_13_io_out ? io_r_398_b : _GEN_5777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5781 = 9'h1 == r_count_14_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5782 = 9'h2 == r_count_14_io_out ? io_r_2_b : _GEN_5781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5783 = 9'h3 == r_count_14_io_out ? io_r_3_b : _GEN_5782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5784 = 9'h4 == r_count_14_io_out ? io_r_4_b : _GEN_5783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5785 = 9'h5 == r_count_14_io_out ? io_r_5_b : _GEN_5784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5786 = 9'h6 == r_count_14_io_out ? io_r_6_b : _GEN_5785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5787 = 9'h7 == r_count_14_io_out ? io_r_7_b : _GEN_5786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5788 = 9'h8 == r_count_14_io_out ? io_r_8_b : _GEN_5787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5789 = 9'h9 == r_count_14_io_out ? io_r_9_b : _GEN_5788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5790 = 9'ha == r_count_14_io_out ? io_r_10_b : _GEN_5789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5791 = 9'hb == r_count_14_io_out ? io_r_11_b : _GEN_5790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5792 = 9'hc == r_count_14_io_out ? io_r_12_b : _GEN_5791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5793 = 9'hd == r_count_14_io_out ? io_r_13_b : _GEN_5792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5794 = 9'he == r_count_14_io_out ? io_r_14_b : _GEN_5793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5795 = 9'hf == r_count_14_io_out ? io_r_15_b : _GEN_5794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5796 = 9'h10 == r_count_14_io_out ? io_r_16_b : _GEN_5795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5797 = 9'h11 == r_count_14_io_out ? io_r_17_b : _GEN_5796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5798 = 9'h12 == r_count_14_io_out ? io_r_18_b : _GEN_5797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5799 = 9'h13 == r_count_14_io_out ? io_r_19_b : _GEN_5798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5800 = 9'h14 == r_count_14_io_out ? io_r_20_b : _GEN_5799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5801 = 9'h15 == r_count_14_io_out ? io_r_21_b : _GEN_5800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5802 = 9'h16 == r_count_14_io_out ? io_r_22_b : _GEN_5801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5803 = 9'h17 == r_count_14_io_out ? io_r_23_b : _GEN_5802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5804 = 9'h18 == r_count_14_io_out ? io_r_24_b : _GEN_5803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5805 = 9'h19 == r_count_14_io_out ? io_r_25_b : _GEN_5804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5806 = 9'h1a == r_count_14_io_out ? io_r_26_b : _GEN_5805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5807 = 9'h1b == r_count_14_io_out ? io_r_27_b : _GEN_5806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5808 = 9'h1c == r_count_14_io_out ? io_r_28_b : _GEN_5807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5809 = 9'h1d == r_count_14_io_out ? io_r_29_b : _GEN_5808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5810 = 9'h1e == r_count_14_io_out ? io_r_30_b : _GEN_5809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5811 = 9'h1f == r_count_14_io_out ? io_r_31_b : _GEN_5810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5812 = 9'h20 == r_count_14_io_out ? io_r_32_b : _GEN_5811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5813 = 9'h21 == r_count_14_io_out ? io_r_33_b : _GEN_5812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5814 = 9'h22 == r_count_14_io_out ? io_r_34_b : _GEN_5813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5815 = 9'h23 == r_count_14_io_out ? io_r_35_b : _GEN_5814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5816 = 9'h24 == r_count_14_io_out ? io_r_36_b : _GEN_5815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5817 = 9'h25 == r_count_14_io_out ? io_r_37_b : _GEN_5816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5818 = 9'h26 == r_count_14_io_out ? io_r_38_b : _GEN_5817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5819 = 9'h27 == r_count_14_io_out ? io_r_39_b : _GEN_5818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5820 = 9'h28 == r_count_14_io_out ? io_r_40_b : _GEN_5819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5821 = 9'h29 == r_count_14_io_out ? io_r_41_b : _GEN_5820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5822 = 9'h2a == r_count_14_io_out ? io_r_42_b : _GEN_5821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5823 = 9'h2b == r_count_14_io_out ? io_r_43_b : _GEN_5822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5824 = 9'h2c == r_count_14_io_out ? io_r_44_b : _GEN_5823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5825 = 9'h2d == r_count_14_io_out ? io_r_45_b : _GEN_5824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5826 = 9'h2e == r_count_14_io_out ? io_r_46_b : _GEN_5825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5827 = 9'h2f == r_count_14_io_out ? io_r_47_b : _GEN_5826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5828 = 9'h30 == r_count_14_io_out ? io_r_48_b : _GEN_5827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5829 = 9'h31 == r_count_14_io_out ? io_r_49_b : _GEN_5828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5830 = 9'h32 == r_count_14_io_out ? io_r_50_b : _GEN_5829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5831 = 9'h33 == r_count_14_io_out ? io_r_51_b : _GEN_5830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5832 = 9'h34 == r_count_14_io_out ? io_r_52_b : _GEN_5831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5833 = 9'h35 == r_count_14_io_out ? io_r_53_b : _GEN_5832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5834 = 9'h36 == r_count_14_io_out ? io_r_54_b : _GEN_5833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5835 = 9'h37 == r_count_14_io_out ? io_r_55_b : _GEN_5834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5836 = 9'h38 == r_count_14_io_out ? io_r_56_b : _GEN_5835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5837 = 9'h39 == r_count_14_io_out ? io_r_57_b : _GEN_5836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5838 = 9'h3a == r_count_14_io_out ? io_r_58_b : _GEN_5837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5839 = 9'h3b == r_count_14_io_out ? io_r_59_b : _GEN_5838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5840 = 9'h3c == r_count_14_io_out ? io_r_60_b : _GEN_5839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5841 = 9'h3d == r_count_14_io_out ? io_r_61_b : _GEN_5840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5842 = 9'h3e == r_count_14_io_out ? io_r_62_b : _GEN_5841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5843 = 9'h3f == r_count_14_io_out ? io_r_63_b : _GEN_5842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5844 = 9'h40 == r_count_14_io_out ? io_r_64_b : _GEN_5843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5845 = 9'h41 == r_count_14_io_out ? io_r_65_b : _GEN_5844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5846 = 9'h42 == r_count_14_io_out ? io_r_66_b : _GEN_5845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5847 = 9'h43 == r_count_14_io_out ? io_r_67_b : _GEN_5846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5848 = 9'h44 == r_count_14_io_out ? io_r_68_b : _GEN_5847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5849 = 9'h45 == r_count_14_io_out ? io_r_69_b : _GEN_5848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5850 = 9'h46 == r_count_14_io_out ? io_r_70_b : _GEN_5849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5851 = 9'h47 == r_count_14_io_out ? io_r_71_b : _GEN_5850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5852 = 9'h48 == r_count_14_io_out ? io_r_72_b : _GEN_5851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5853 = 9'h49 == r_count_14_io_out ? io_r_73_b : _GEN_5852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5854 = 9'h4a == r_count_14_io_out ? io_r_74_b : _GEN_5853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5855 = 9'h4b == r_count_14_io_out ? io_r_75_b : _GEN_5854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5856 = 9'h4c == r_count_14_io_out ? io_r_76_b : _GEN_5855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5857 = 9'h4d == r_count_14_io_out ? io_r_77_b : _GEN_5856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5858 = 9'h4e == r_count_14_io_out ? io_r_78_b : _GEN_5857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5859 = 9'h4f == r_count_14_io_out ? io_r_79_b : _GEN_5858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5860 = 9'h50 == r_count_14_io_out ? io_r_80_b : _GEN_5859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5861 = 9'h51 == r_count_14_io_out ? io_r_81_b : _GEN_5860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5862 = 9'h52 == r_count_14_io_out ? io_r_82_b : _GEN_5861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5863 = 9'h53 == r_count_14_io_out ? io_r_83_b : _GEN_5862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5864 = 9'h54 == r_count_14_io_out ? io_r_84_b : _GEN_5863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5865 = 9'h55 == r_count_14_io_out ? io_r_85_b : _GEN_5864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5866 = 9'h56 == r_count_14_io_out ? io_r_86_b : _GEN_5865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5867 = 9'h57 == r_count_14_io_out ? io_r_87_b : _GEN_5866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5868 = 9'h58 == r_count_14_io_out ? io_r_88_b : _GEN_5867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5869 = 9'h59 == r_count_14_io_out ? io_r_89_b : _GEN_5868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5870 = 9'h5a == r_count_14_io_out ? io_r_90_b : _GEN_5869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5871 = 9'h5b == r_count_14_io_out ? io_r_91_b : _GEN_5870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5872 = 9'h5c == r_count_14_io_out ? io_r_92_b : _GEN_5871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5873 = 9'h5d == r_count_14_io_out ? io_r_93_b : _GEN_5872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5874 = 9'h5e == r_count_14_io_out ? io_r_94_b : _GEN_5873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5875 = 9'h5f == r_count_14_io_out ? io_r_95_b : _GEN_5874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5876 = 9'h60 == r_count_14_io_out ? io_r_96_b : _GEN_5875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5877 = 9'h61 == r_count_14_io_out ? io_r_97_b : _GEN_5876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5878 = 9'h62 == r_count_14_io_out ? io_r_98_b : _GEN_5877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5879 = 9'h63 == r_count_14_io_out ? io_r_99_b : _GEN_5878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5880 = 9'h64 == r_count_14_io_out ? io_r_100_b : _GEN_5879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5881 = 9'h65 == r_count_14_io_out ? io_r_101_b : _GEN_5880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5882 = 9'h66 == r_count_14_io_out ? io_r_102_b : _GEN_5881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5883 = 9'h67 == r_count_14_io_out ? io_r_103_b : _GEN_5882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5884 = 9'h68 == r_count_14_io_out ? io_r_104_b : _GEN_5883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5885 = 9'h69 == r_count_14_io_out ? io_r_105_b : _GEN_5884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5886 = 9'h6a == r_count_14_io_out ? io_r_106_b : _GEN_5885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5887 = 9'h6b == r_count_14_io_out ? io_r_107_b : _GEN_5886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5888 = 9'h6c == r_count_14_io_out ? io_r_108_b : _GEN_5887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5889 = 9'h6d == r_count_14_io_out ? io_r_109_b : _GEN_5888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5890 = 9'h6e == r_count_14_io_out ? io_r_110_b : _GEN_5889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5891 = 9'h6f == r_count_14_io_out ? io_r_111_b : _GEN_5890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5892 = 9'h70 == r_count_14_io_out ? io_r_112_b : _GEN_5891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5893 = 9'h71 == r_count_14_io_out ? io_r_113_b : _GEN_5892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5894 = 9'h72 == r_count_14_io_out ? io_r_114_b : _GEN_5893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5895 = 9'h73 == r_count_14_io_out ? io_r_115_b : _GEN_5894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5896 = 9'h74 == r_count_14_io_out ? io_r_116_b : _GEN_5895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5897 = 9'h75 == r_count_14_io_out ? io_r_117_b : _GEN_5896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5898 = 9'h76 == r_count_14_io_out ? io_r_118_b : _GEN_5897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5899 = 9'h77 == r_count_14_io_out ? io_r_119_b : _GEN_5898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5900 = 9'h78 == r_count_14_io_out ? io_r_120_b : _GEN_5899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5901 = 9'h79 == r_count_14_io_out ? io_r_121_b : _GEN_5900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5902 = 9'h7a == r_count_14_io_out ? io_r_122_b : _GEN_5901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5903 = 9'h7b == r_count_14_io_out ? io_r_123_b : _GEN_5902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5904 = 9'h7c == r_count_14_io_out ? io_r_124_b : _GEN_5903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5905 = 9'h7d == r_count_14_io_out ? io_r_125_b : _GEN_5904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5906 = 9'h7e == r_count_14_io_out ? io_r_126_b : _GEN_5905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5907 = 9'h7f == r_count_14_io_out ? io_r_127_b : _GEN_5906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5908 = 9'h80 == r_count_14_io_out ? io_r_128_b : _GEN_5907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5909 = 9'h81 == r_count_14_io_out ? io_r_129_b : _GEN_5908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5910 = 9'h82 == r_count_14_io_out ? io_r_130_b : _GEN_5909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5911 = 9'h83 == r_count_14_io_out ? io_r_131_b : _GEN_5910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5912 = 9'h84 == r_count_14_io_out ? io_r_132_b : _GEN_5911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5913 = 9'h85 == r_count_14_io_out ? io_r_133_b : _GEN_5912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5914 = 9'h86 == r_count_14_io_out ? io_r_134_b : _GEN_5913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5915 = 9'h87 == r_count_14_io_out ? io_r_135_b : _GEN_5914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5916 = 9'h88 == r_count_14_io_out ? io_r_136_b : _GEN_5915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5917 = 9'h89 == r_count_14_io_out ? io_r_137_b : _GEN_5916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5918 = 9'h8a == r_count_14_io_out ? io_r_138_b : _GEN_5917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5919 = 9'h8b == r_count_14_io_out ? io_r_139_b : _GEN_5918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5920 = 9'h8c == r_count_14_io_out ? io_r_140_b : _GEN_5919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5921 = 9'h8d == r_count_14_io_out ? io_r_141_b : _GEN_5920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5922 = 9'h8e == r_count_14_io_out ? io_r_142_b : _GEN_5921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5923 = 9'h8f == r_count_14_io_out ? io_r_143_b : _GEN_5922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5924 = 9'h90 == r_count_14_io_out ? io_r_144_b : _GEN_5923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5925 = 9'h91 == r_count_14_io_out ? io_r_145_b : _GEN_5924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5926 = 9'h92 == r_count_14_io_out ? io_r_146_b : _GEN_5925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5927 = 9'h93 == r_count_14_io_out ? io_r_147_b : _GEN_5926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5928 = 9'h94 == r_count_14_io_out ? io_r_148_b : _GEN_5927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5929 = 9'h95 == r_count_14_io_out ? io_r_149_b : _GEN_5928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5930 = 9'h96 == r_count_14_io_out ? io_r_150_b : _GEN_5929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5931 = 9'h97 == r_count_14_io_out ? io_r_151_b : _GEN_5930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5932 = 9'h98 == r_count_14_io_out ? io_r_152_b : _GEN_5931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5933 = 9'h99 == r_count_14_io_out ? io_r_153_b : _GEN_5932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5934 = 9'h9a == r_count_14_io_out ? io_r_154_b : _GEN_5933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5935 = 9'h9b == r_count_14_io_out ? io_r_155_b : _GEN_5934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5936 = 9'h9c == r_count_14_io_out ? io_r_156_b : _GEN_5935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5937 = 9'h9d == r_count_14_io_out ? io_r_157_b : _GEN_5936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5938 = 9'h9e == r_count_14_io_out ? io_r_158_b : _GEN_5937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5939 = 9'h9f == r_count_14_io_out ? io_r_159_b : _GEN_5938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5940 = 9'ha0 == r_count_14_io_out ? io_r_160_b : _GEN_5939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5941 = 9'ha1 == r_count_14_io_out ? io_r_161_b : _GEN_5940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5942 = 9'ha2 == r_count_14_io_out ? io_r_162_b : _GEN_5941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5943 = 9'ha3 == r_count_14_io_out ? io_r_163_b : _GEN_5942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5944 = 9'ha4 == r_count_14_io_out ? io_r_164_b : _GEN_5943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5945 = 9'ha5 == r_count_14_io_out ? io_r_165_b : _GEN_5944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5946 = 9'ha6 == r_count_14_io_out ? io_r_166_b : _GEN_5945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5947 = 9'ha7 == r_count_14_io_out ? io_r_167_b : _GEN_5946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5948 = 9'ha8 == r_count_14_io_out ? io_r_168_b : _GEN_5947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5949 = 9'ha9 == r_count_14_io_out ? io_r_169_b : _GEN_5948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5950 = 9'haa == r_count_14_io_out ? io_r_170_b : _GEN_5949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5951 = 9'hab == r_count_14_io_out ? io_r_171_b : _GEN_5950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5952 = 9'hac == r_count_14_io_out ? io_r_172_b : _GEN_5951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5953 = 9'had == r_count_14_io_out ? io_r_173_b : _GEN_5952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5954 = 9'hae == r_count_14_io_out ? io_r_174_b : _GEN_5953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5955 = 9'haf == r_count_14_io_out ? io_r_175_b : _GEN_5954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5956 = 9'hb0 == r_count_14_io_out ? io_r_176_b : _GEN_5955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5957 = 9'hb1 == r_count_14_io_out ? io_r_177_b : _GEN_5956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5958 = 9'hb2 == r_count_14_io_out ? io_r_178_b : _GEN_5957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5959 = 9'hb3 == r_count_14_io_out ? io_r_179_b : _GEN_5958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5960 = 9'hb4 == r_count_14_io_out ? io_r_180_b : _GEN_5959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5961 = 9'hb5 == r_count_14_io_out ? io_r_181_b : _GEN_5960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5962 = 9'hb6 == r_count_14_io_out ? io_r_182_b : _GEN_5961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5963 = 9'hb7 == r_count_14_io_out ? io_r_183_b : _GEN_5962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5964 = 9'hb8 == r_count_14_io_out ? io_r_184_b : _GEN_5963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5965 = 9'hb9 == r_count_14_io_out ? io_r_185_b : _GEN_5964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5966 = 9'hba == r_count_14_io_out ? io_r_186_b : _GEN_5965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5967 = 9'hbb == r_count_14_io_out ? io_r_187_b : _GEN_5966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5968 = 9'hbc == r_count_14_io_out ? io_r_188_b : _GEN_5967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5969 = 9'hbd == r_count_14_io_out ? io_r_189_b : _GEN_5968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5970 = 9'hbe == r_count_14_io_out ? io_r_190_b : _GEN_5969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5971 = 9'hbf == r_count_14_io_out ? io_r_191_b : _GEN_5970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5972 = 9'hc0 == r_count_14_io_out ? io_r_192_b : _GEN_5971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5973 = 9'hc1 == r_count_14_io_out ? io_r_193_b : _GEN_5972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5974 = 9'hc2 == r_count_14_io_out ? io_r_194_b : _GEN_5973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5975 = 9'hc3 == r_count_14_io_out ? io_r_195_b : _GEN_5974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5976 = 9'hc4 == r_count_14_io_out ? io_r_196_b : _GEN_5975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5977 = 9'hc5 == r_count_14_io_out ? io_r_197_b : _GEN_5976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5978 = 9'hc6 == r_count_14_io_out ? io_r_198_b : _GEN_5977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5979 = 9'hc7 == r_count_14_io_out ? io_r_199_b : _GEN_5978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5980 = 9'hc8 == r_count_14_io_out ? io_r_200_b : _GEN_5979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5981 = 9'hc9 == r_count_14_io_out ? io_r_201_b : _GEN_5980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5982 = 9'hca == r_count_14_io_out ? io_r_202_b : _GEN_5981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5983 = 9'hcb == r_count_14_io_out ? io_r_203_b : _GEN_5982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5984 = 9'hcc == r_count_14_io_out ? io_r_204_b : _GEN_5983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5985 = 9'hcd == r_count_14_io_out ? io_r_205_b : _GEN_5984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5986 = 9'hce == r_count_14_io_out ? io_r_206_b : _GEN_5985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5987 = 9'hcf == r_count_14_io_out ? io_r_207_b : _GEN_5986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5988 = 9'hd0 == r_count_14_io_out ? io_r_208_b : _GEN_5987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5989 = 9'hd1 == r_count_14_io_out ? io_r_209_b : _GEN_5988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5990 = 9'hd2 == r_count_14_io_out ? io_r_210_b : _GEN_5989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5991 = 9'hd3 == r_count_14_io_out ? io_r_211_b : _GEN_5990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5992 = 9'hd4 == r_count_14_io_out ? io_r_212_b : _GEN_5991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5993 = 9'hd5 == r_count_14_io_out ? io_r_213_b : _GEN_5992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5994 = 9'hd6 == r_count_14_io_out ? io_r_214_b : _GEN_5993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5995 = 9'hd7 == r_count_14_io_out ? io_r_215_b : _GEN_5994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5996 = 9'hd8 == r_count_14_io_out ? io_r_216_b : _GEN_5995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5997 = 9'hd9 == r_count_14_io_out ? io_r_217_b : _GEN_5996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5998 = 9'hda == r_count_14_io_out ? io_r_218_b : _GEN_5997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5999 = 9'hdb == r_count_14_io_out ? io_r_219_b : _GEN_5998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6000 = 9'hdc == r_count_14_io_out ? io_r_220_b : _GEN_5999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6001 = 9'hdd == r_count_14_io_out ? io_r_221_b : _GEN_6000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6002 = 9'hde == r_count_14_io_out ? io_r_222_b : _GEN_6001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6003 = 9'hdf == r_count_14_io_out ? io_r_223_b : _GEN_6002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6004 = 9'he0 == r_count_14_io_out ? io_r_224_b : _GEN_6003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6005 = 9'he1 == r_count_14_io_out ? io_r_225_b : _GEN_6004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6006 = 9'he2 == r_count_14_io_out ? io_r_226_b : _GEN_6005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6007 = 9'he3 == r_count_14_io_out ? io_r_227_b : _GEN_6006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6008 = 9'he4 == r_count_14_io_out ? io_r_228_b : _GEN_6007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6009 = 9'he5 == r_count_14_io_out ? io_r_229_b : _GEN_6008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6010 = 9'he6 == r_count_14_io_out ? io_r_230_b : _GEN_6009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6011 = 9'he7 == r_count_14_io_out ? io_r_231_b : _GEN_6010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6012 = 9'he8 == r_count_14_io_out ? io_r_232_b : _GEN_6011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6013 = 9'he9 == r_count_14_io_out ? io_r_233_b : _GEN_6012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6014 = 9'hea == r_count_14_io_out ? io_r_234_b : _GEN_6013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6015 = 9'heb == r_count_14_io_out ? io_r_235_b : _GEN_6014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6016 = 9'hec == r_count_14_io_out ? io_r_236_b : _GEN_6015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6017 = 9'hed == r_count_14_io_out ? io_r_237_b : _GEN_6016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6018 = 9'hee == r_count_14_io_out ? io_r_238_b : _GEN_6017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6019 = 9'hef == r_count_14_io_out ? io_r_239_b : _GEN_6018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6020 = 9'hf0 == r_count_14_io_out ? io_r_240_b : _GEN_6019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6021 = 9'hf1 == r_count_14_io_out ? io_r_241_b : _GEN_6020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6022 = 9'hf2 == r_count_14_io_out ? io_r_242_b : _GEN_6021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6023 = 9'hf3 == r_count_14_io_out ? io_r_243_b : _GEN_6022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6024 = 9'hf4 == r_count_14_io_out ? io_r_244_b : _GEN_6023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6025 = 9'hf5 == r_count_14_io_out ? io_r_245_b : _GEN_6024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6026 = 9'hf6 == r_count_14_io_out ? io_r_246_b : _GEN_6025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6027 = 9'hf7 == r_count_14_io_out ? io_r_247_b : _GEN_6026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6028 = 9'hf8 == r_count_14_io_out ? io_r_248_b : _GEN_6027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6029 = 9'hf9 == r_count_14_io_out ? io_r_249_b : _GEN_6028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6030 = 9'hfa == r_count_14_io_out ? io_r_250_b : _GEN_6029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6031 = 9'hfb == r_count_14_io_out ? io_r_251_b : _GEN_6030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6032 = 9'hfc == r_count_14_io_out ? io_r_252_b : _GEN_6031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6033 = 9'hfd == r_count_14_io_out ? io_r_253_b : _GEN_6032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6034 = 9'hfe == r_count_14_io_out ? io_r_254_b : _GEN_6033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6035 = 9'hff == r_count_14_io_out ? io_r_255_b : _GEN_6034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6036 = 9'h100 == r_count_14_io_out ? io_r_256_b : _GEN_6035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6037 = 9'h101 == r_count_14_io_out ? io_r_257_b : _GEN_6036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6038 = 9'h102 == r_count_14_io_out ? io_r_258_b : _GEN_6037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6039 = 9'h103 == r_count_14_io_out ? io_r_259_b : _GEN_6038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6040 = 9'h104 == r_count_14_io_out ? io_r_260_b : _GEN_6039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6041 = 9'h105 == r_count_14_io_out ? io_r_261_b : _GEN_6040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6042 = 9'h106 == r_count_14_io_out ? io_r_262_b : _GEN_6041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6043 = 9'h107 == r_count_14_io_out ? io_r_263_b : _GEN_6042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6044 = 9'h108 == r_count_14_io_out ? io_r_264_b : _GEN_6043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6045 = 9'h109 == r_count_14_io_out ? io_r_265_b : _GEN_6044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6046 = 9'h10a == r_count_14_io_out ? io_r_266_b : _GEN_6045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6047 = 9'h10b == r_count_14_io_out ? io_r_267_b : _GEN_6046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6048 = 9'h10c == r_count_14_io_out ? io_r_268_b : _GEN_6047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6049 = 9'h10d == r_count_14_io_out ? io_r_269_b : _GEN_6048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6050 = 9'h10e == r_count_14_io_out ? io_r_270_b : _GEN_6049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6051 = 9'h10f == r_count_14_io_out ? io_r_271_b : _GEN_6050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6052 = 9'h110 == r_count_14_io_out ? io_r_272_b : _GEN_6051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6053 = 9'h111 == r_count_14_io_out ? io_r_273_b : _GEN_6052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6054 = 9'h112 == r_count_14_io_out ? io_r_274_b : _GEN_6053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6055 = 9'h113 == r_count_14_io_out ? io_r_275_b : _GEN_6054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6056 = 9'h114 == r_count_14_io_out ? io_r_276_b : _GEN_6055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6057 = 9'h115 == r_count_14_io_out ? io_r_277_b : _GEN_6056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6058 = 9'h116 == r_count_14_io_out ? io_r_278_b : _GEN_6057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6059 = 9'h117 == r_count_14_io_out ? io_r_279_b : _GEN_6058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6060 = 9'h118 == r_count_14_io_out ? io_r_280_b : _GEN_6059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6061 = 9'h119 == r_count_14_io_out ? io_r_281_b : _GEN_6060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6062 = 9'h11a == r_count_14_io_out ? io_r_282_b : _GEN_6061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6063 = 9'h11b == r_count_14_io_out ? io_r_283_b : _GEN_6062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6064 = 9'h11c == r_count_14_io_out ? io_r_284_b : _GEN_6063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6065 = 9'h11d == r_count_14_io_out ? io_r_285_b : _GEN_6064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6066 = 9'h11e == r_count_14_io_out ? io_r_286_b : _GEN_6065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6067 = 9'h11f == r_count_14_io_out ? io_r_287_b : _GEN_6066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6068 = 9'h120 == r_count_14_io_out ? io_r_288_b : _GEN_6067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6069 = 9'h121 == r_count_14_io_out ? io_r_289_b : _GEN_6068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6070 = 9'h122 == r_count_14_io_out ? io_r_290_b : _GEN_6069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6071 = 9'h123 == r_count_14_io_out ? io_r_291_b : _GEN_6070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6072 = 9'h124 == r_count_14_io_out ? io_r_292_b : _GEN_6071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6073 = 9'h125 == r_count_14_io_out ? io_r_293_b : _GEN_6072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6074 = 9'h126 == r_count_14_io_out ? io_r_294_b : _GEN_6073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6075 = 9'h127 == r_count_14_io_out ? io_r_295_b : _GEN_6074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6076 = 9'h128 == r_count_14_io_out ? io_r_296_b : _GEN_6075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6077 = 9'h129 == r_count_14_io_out ? io_r_297_b : _GEN_6076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6078 = 9'h12a == r_count_14_io_out ? io_r_298_b : _GEN_6077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6079 = 9'h12b == r_count_14_io_out ? io_r_299_b : _GEN_6078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6080 = 9'h12c == r_count_14_io_out ? io_r_300_b : _GEN_6079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6081 = 9'h12d == r_count_14_io_out ? io_r_301_b : _GEN_6080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6082 = 9'h12e == r_count_14_io_out ? io_r_302_b : _GEN_6081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6083 = 9'h12f == r_count_14_io_out ? io_r_303_b : _GEN_6082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6084 = 9'h130 == r_count_14_io_out ? io_r_304_b : _GEN_6083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6085 = 9'h131 == r_count_14_io_out ? io_r_305_b : _GEN_6084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6086 = 9'h132 == r_count_14_io_out ? io_r_306_b : _GEN_6085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6087 = 9'h133 == r_count_14_io_out ? io_r_307_b : _GEN_6086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6088 = 9'h134 == r_count_14_io_out ? io_r_308_b : _GEN_6087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6089 = 9'h135 == r_count_14_io_out ? io_r_309_b : _GEN_6088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6090 = 9'h136 == r_count_14_io_out ? io_r_310_b : _GEN_6089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6091 = 9'h137 == r_count_14_io_out ? io_r_311_b : _GEN_6090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6092 = 9'h138 == r_count_14_io_out ? io_r_312_b : _GEN_6091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6093 = 9'h139 == r_count_14_io_out ? io_r_313_b : _GEN_6092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6094 = 9'h13a == r_count_14_io_out ? io_r_314_b : _GEN_6093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6095 = 9'h13b == r_count_14_io_out ? io_r_315_b : _GEN_6094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6096 = 9'h13c == r_count_14_io_out ? io_r_316_b : _GEN_6095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6097 = 9'h13d == r_count_14_io_out ? io_r_317_b : _GEN_6096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6098 = 9'h13e == r_count_14_io_out ? io_r_318_b : _GEN_6097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6099 = 9'h13f == r_count_14_io_out ? io_r_319_b : _GEN_6098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6100 = 9'h140 == r_count_14_io_out ? io_r_320_b : _GEN_6099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6101 = 9'h141 == r_count_14_io_out ? io_r_321_b : _GEN_6100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6102 = 9'h142 == r_count_14_io_out ? io_r_322_b : _GEN_6101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6103 = 9'h143 == r_count_14_io_out ? io_r_323_b : _GEN_6102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6104 = 9'h144 == r_count_14_io_out ? io_r_324_b : _GEN_6103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6105 = 9'h145 == r_count_14_io_out ? io_r_325_b : _GEN_6104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6106 = 9'h146 == r_count_14_io_out ? io_r_326_b : _GEN_6105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6107 = 9'h147 == r_count_14_io_out ? io_r_327_b : _GEN_6106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6108 = 9'h148 == r_count_14_io_out ? io_r_328_b : _GEN_6107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6109 = 9'h149 == r_count_14_io_out ? io_r_329_b : _GEN_6108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6110 = 9'h14a == r_count_14_io_out ? io_r_330_b : _GEN_6109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6111 = 9'h14b == r_count_14_io_out ? io_r_331_b : _GEN_6110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6112 = 9'h14c == r_count_14_io_out ? io_r_332_b : _GEN_6111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6113 = 9'h14d == r_count_14_io_out ? io_r_333_b : _GEN_6112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6114 = 9'h14e == r_count_14_io_out ? io_r_334_b : _GEN_6113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6115 = 9'h14f == r_count_14_io_out ? io_r_335_b : _GEN_6114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6116 = 9'h150 == r_count_14_io_out ? io_r_336_b : _GEN_6115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6117 = 9'h151 == r_count_14_io_out ? io_r_337_b : _GEN_6116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6118 = 9'h152 == r_count_14_io_out ? io_r_338_b : _GEN_6117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6119 = 9'h153 == r_count_14_io_out ? io_r_339_b : _GEN_6118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6120 = 9'h154 == r_count_14_io_out ? io_r_340_b : _GEN_6119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6121 = 9'h155 == r_count_14_io_out ? io_r_341_b : _GEN_6120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6122 = 9'h156 == r_count_14_io_out ? io_r_342_b : _GEN_6121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6123 = 9'h157 == r_count_14_io_out ? io_r_343_b : _GEN_6122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6124 = 9'h158 == r_count_14_io_out ? io_r_344_b : _GEN_6123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6125 = 9'h159 == r_count_14_io_out ? io_r_345_b : _GEN_6124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6126 = 9'h15a == r_count_14_io_out ? io_r_346_b : _GEN_6125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6127 = 9'h15b == r_count_14_io_out ? io_r_347_b : _GEN_6126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6128 = 9'h15c == r_count_14_io_out ? io_r_348_b : _GEN_6127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6129 = 9'h15d == r_count_14_io_out ? io_r_349_b : _GEN_6128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6130 = 9'h15e == r_count_14_io_out ? io_r_350_b : _GEN_6129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6131 = 9'h15f == r_count_14_io_out ? io_r_351_b : _GEN_6130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6132 = 9'h160 == r_count_14_io_out ? io_r_352_b : _GEN_6131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6133 = 9'h161 == r_count_14_io_out ? io_r_353_b : _GEN_6132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6134 = 9'h162 == r_count_14_io_out ? io_r_354_b : _GEN_6133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6135 = 9'h163 == r_count_14_io_out ? io_r_355_b : _GEN_6134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6136 = 9'h164 == r_count_14_io_out ? io_r_356_b : _GEN_6135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6137 = 9'h165 == r_count_14_io_out ? io_r_357_b : _GEN_6136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6138 = 9'h166 == r_count_14_io_out ? io_r_358_b : _GEN_6137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6139 = 9'h167 == r_count_14_io_out ? io_r_359_b : _GEN_6138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6140 = 9'h168 == r_count_14_io_out ? io_r_360_b : _GEN_6139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6141 = 9'h169 == r_count_14_io_out ? io_r_361_b : _GEN_6140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6142 = 9'h16a == r_count_14_io_out ? io_r_362_b : _GEN_6141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6143 = 9'h16b == r_count_14_io_out ? io_r_363_b : _GEN_6142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6144 = 9'h16c == r_count_14_io_out ? io_r_364_b : _GEN_6143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6145 = 9'h16d == r_count_14_io_out ? io_r_365_b : _GEN_6144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6146 = 9'h16e == r_count_14_io_out ? io_r_366_b : _GEN_6145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6147 = 9'h16f == r_count_14_io_out ? io_r_367_b : _GEN_6146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6148 = 9'h170 == r_count_14_io_out ? io_r_368_b : _GEN_6147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6149 = 9'h171 == r_count_14_io_out ? io_r_369_b : _GEN_6148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6150 = 9'h172 == r_count_14_io_out ? io_r_370_b : _GEN_6149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6151 = 9'h173 == r_count_14_io_out ? io_r_371_b : _GEN_6150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6152 = 9'h174 == r_count_14_io_out ? io_r_372_b : _GEN_6151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6153 = 9'h175 == r_count_14_io_out ? io_r_373_b : _GEN_6152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6154 = 9'h176 == r_count_14_io_out ? io_r_374_b : _GEN_6153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6155 = 9'h177 == r_count_14_io_out ? io_r_375_b : _GEN_6154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6156 = 9'h178 == r_count_14_io_out ? io_r_376_b : _GEN_6155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6157 = 9'h179 == r_count_14_io_out ? io_r_377_b : _GEN_6156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6158 = 9'h17a == r_count_14_io_out ? io_r_378_b : _GEN_6157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6159 = 9'h17b == r_count_14_io_out ? io_r_379_b : _GEN_6158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6160 = 9'h17c == r_count_14_io_out ? io_r_380_b : _GEN_6159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6161 = 9'h17d == r_count_14_io_out ? io_r_381_b : _GEN_6160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6162 = 9'h17e == r_count_14_io_out ? io_r_382_b : _GEN_6161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6163 = 9'h17f == r_count_14_io_out ? io_r_383_b : _GEN_6162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6164 = 9'h180 == r_count_14_io_out ? io_r_384_b : _GEN_6163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6165 = 9'h181 == r_count_14_io_out ? io_r_385_b : _GEN_6164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6166 = 9'h182 == r_count_14_io_out ? io_r_386_b : _GEN_6165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6167 = 9'h183 == r_count_14_io_out ? io_r_387_b : _GEN_6166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6168 = 9'h184 == r_count_14_io_out ? io_r_388_b : _GEN_6167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6169 = 9'h185 == r_count_14_io_out ? io_r_389_b : _GEN_6168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6170 = 9'h186 == r_count_14_io_out ? io_r_390_b : _GEN_6169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6171 = 9'h187 == r_count_14_io_out ? io_r_391_b : _GEN_6170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6172 = 9'h188 == r_count_14_io_out ? io_r_392_b : _GEN_6171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6173 = 9'h189 == r_count_14_io_out ? io_r_393_b : _GEN_6172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6174 = 9'h18a == r_count_14_io_out ? io_r_394_b : _GEN_6173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6175 = 9'h18b == r_count_14_io_out ? io_r_395_b : _GEN_6174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6176 = 9'h18c == r_count_14_io_out ? io_r_396_b : _GEN_6175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6177 = 9'h18d == r_count_14_io_out ? io_r_397_b : _GEN_6176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6178 = 9'h18e == r_count_14_io_out ? io_r_398_b : _GEN_6177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6181 = 9'h1 == r_count_15_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6182 = 9'h2 == r_count_15_io_out ? io_r_2_b : _GEN_6181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6183 = 9'h3 == r_count_15_io_out ? io_r_3_b : _GEN_6182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6184 = 9'h4 == r_count_15_io_out ? io_r_4_b : _GEN_6183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6185 = 9'h5 == r_count_15_io_out ? io_r_5_b : _GEN_6184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6186 = 9'h6 == r_count_15_io_out ? io_r_6_b : _GEN_6185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6187 = 9'h7 == r_count_15_io_out ? io_r_7_b : _GEN_6186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6188 = 9'h8 == r_count_15_io_out ? io_r_8_b : _GEN_6187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6189 = 9'h9 == r_count_15_io_out ? io_r_9_b : _GEN_6188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6190 = 9'ha == r_count_15_io_out ? io_r_10_b : _GEN_6189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6191 = 9'hb == r_count_15_io_out ? io_r_11_b : _GEN_6190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6192 = 9'hc == r_count_15_io_out ? io_r_12_b : _GEN_6191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6193 = 9'hd == r_count_15_io_out ? io_r_13_b : _GEN_6192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6194 = 9'he == r_count_15_io_out ? io_r_14_b : _GEN_6193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6195 = 9'hf == r_count_15_io_out ? io_r_15_b : _GEN_6194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6196 = 9'h10 == r_count_15_io_out ? io_r_16_b : _GEN_6195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6197 = 9'h11 == r_count_15_io_out ? io_r_17_b : _GEN_6196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6198 = 9'h12 == r_count_15_io_out ? io_r_18_b : _GEN_6197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6199 = 9'h13 == r_count_15_io_out ? io_r_19_b : _GEN_6198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6200 = 9'h14 == r_count_15_io_out ? io_r_20_b : _GEN_6199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6201 = 9'h15 == r_count_15_io_out ? io_r_21_b : _GEN_6200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6202 = 9'h16 == r_count_15_io_out ? io_r_22_b : _GEN_6201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6203 = 9'h17 == r_count_15_io_out ? io_r_23_b : _GEN_6202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6204 = 9'h18 == r_count_15_io_out ? io_r_24_b : _GEN_6203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6205 = 9'h19 == r_count_15_io_out ? io_r_25_b : _GEN_6204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6206 = 9'h1a == r_count_15_io_out ? io_r_26_b : _GEN_6205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6207 = 9'h1b == r_count_15_io_out ? io_r_27_b : _GEN_6206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6208 = 9'h1c == r_count_15_io_out ? io_r_28_b : _GEN_6207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6209 = 9'h1d == r_count_15_io_out ? io_r_29_b : _GEN_6208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6210 = 9'h1e == r_count_15_io_out ? io_r_30_b : _GEN_6209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6211 = 9'h1f == r_count_15_io_out ? io_r_31_b : _GEN_6210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6212 = 9'h20 == r_count_15_io_out ? io_r_32_b : _GEN_6211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6213 = 9'h21 == r_count_15_io_out ? io_r_33_b : _GEN_6212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6214 = 9'h22 == r_count_15_io_out ? io_r_34_b : _GEN_6213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6215 = 9'h23 == r_count_15_io_out ? io_r_35_b : _GEN_6214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6216 = 9'h24 == r_count_15_io_out ? io_r_36_b : _GEN_6215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6217 = 9'h25 == r_count_15_io_out ? io_r_37_b : _GEN_6216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6218 = 9'h26 == r_count_15_io_out ? io_r_38_b : _GEN_6217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6219 = 9'h27 == r_count_15_io_out ? io_r_39_b : _GEN_6218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6220 = 9'h28 == r_count_15_io_out ? io_r_40_b : _GEN_6219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6221 = 9'h29 == r_count_15_io_out ? io_r_41_b : _GEN_6220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6222 = 9'h2a == r_count_15_io_out ? io_r_42_b : _GEN_6221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6223 = 9'h2b == r_count_15_io_out ? io_r_43_b : _GEN_6222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6224 = 9'h2c == r_count_15_io_out ? io_r_44_b : _GEN_6223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6225 = 9'h2d == r_count_15_io_out ? io_r_45_b : _GEN_6224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6226 = 9'h2e == r_count_15_io_out ? io_r_46_b : _GEN_6225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6227 = 9'h2f == r_count_15_io_out ? io_r_47_b : _GEN_6226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6228 = 9'h30 == r_count_15_io_out ? io_r_48_b : _GEN_6227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6229 = 9'h31 == r_count_15_io_out ? io_r_49_b : _GEN_6228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6230 = 9'h32 == r_count_15_io_out ? io_r_50_b : _GEN_6229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6231 = 9'h33 == r_count_15_io_out ? io_r_51_b : _GEN_6230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6232 = 9'h34 == r_count_15_io_out ? io_r_52_b : _GEN_6231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6233 = 9'h35 == r_count_15_io_out ? io_r_53_b : _GEN_6232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6234 = 9'h36 == r_count_15_io_out ? io_r_54_b : _GEN_6233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6235 = 9'h37 == r_count_15_io_out ? io_r_55_b : _GEN_6234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6236 = 9'h38 == r_count_15_io_out ? io_r_56_b : _GEN_6235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6237 = 9'h39 == r_count_15_io_out ? io_r_57_b : _GEN_6236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6238 = 9'h3a == r_count_15_io_out ? io_r_58_b : _GEN_6237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6239 = 9'h3b == r_count_15_io_out ? io_r_59_b : _GEN_6238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6240 = 9'h3c == r_count_15_io_out ? io_r_60_b : _GEN_6239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6241 = 9'h3d == r_count_15_io_out ? io_r_61_b : _GEN_6240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6242 = 9'h3e == r_count_15_io_out ? io_r_62_b : _GEN_6241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6243 = 9'h3f == r_count_15_io_out ? io_r_63_b : _GEN_6242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6244 = 9'h40 == r_count_15_io_out ? io_r_64_b : _GEN_6243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6245 = 9'h41 == r_count_15_io_out ? io_r_65_b : _GEN_6244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6246 = 9'h42 == r_count_15_io_out ? io_r_66_b : _GEN_6245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6247 = 9'h43 == r_count_15_io_out ? io_r_67_b : _GEN_6246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6248 = 9'h44 == r_count_15_io_out ? io_r_68_b : _GEN_6247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6249 = 9'h45 == r_count_15_io_out ? io_r_69_b : _GEN_6248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6250 = 9'h46 == r_count_15_io_out ? io_r_70_b : _GEN_6249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6251 = 9'h47 == r_count_15_io_out ? io_r_71_b : _GEN_6250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6252 = 9'h48 == r_count_15_io_out ? io_r_72_b : _GEN_6251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6253 = 9'h49 == r_count_15_io_out ? io_r_73_b : _GEN_6252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6254 = 9'h4a == r_count_15_io_out ? io_r_74_b : _GEN_6253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6255 = 9'h4b == r_count_15_io_out ? io_r_75_b : _GEN_6254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6256 = 9'h4c == r_count_15_io_out ? io_r_76_b : _GEN_6255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6257 = 9'h4d == r_count_15_io_out ? io_r_77_b : _GEN_6256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6258 = 9'h4e == r_count_15_io_out ? io_r_78_b : _GEN_6257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6259 = 9'h4f == r_count_15_io_out ? io_r_79_b : _GEN_6258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6260 = 9'h50 == r_count_15_io_out ? io_r_80_b : _GEN_6259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6261 = 9'h51 == r_count_15_io_out ? io_r_81_b : _GEN_6260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6262 = 9'h52 == r_count_15_io_out ? io_r_82_b : _GEN_6261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6263 = 9'h53 == r_count_15_io_out ? io_r_83_b : _GEN_6262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6264 = 9'h54 == r_count_15_io_out ? io_r_84_b : _GEN_6263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6265 = 9'h55 == r_count_15_io_out ? io_r_85_b : _GEN_6264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6266 = 9'h56 == r_count_15_io_out ? io_r_86_b : _GEN_6265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6267 = 9'h57 == r_count_15_io_out ? io_r_87_b : _GEN_6266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6268 = 9'h58 == r_count_15_io_out ? io_r_88_b : _GEN_6267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6269 = 9'h59 == r_count_15_io_out ? io_r_89_b : _GEN_6268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6270 = 9'h5a == r_count_15_io_out ? io_r_90_b : _GEN_6269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6271 = 9'h5b == r_count_15_io_out ? io_r_91_b : _GEN_6270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6272 = 9'h5c == r_count_15_io_out ? io_r_92_b : _GEN_6271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6273 = 9'h5d == r_count_15_io_out ? io_r_93_b : _GEN_6272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6274 = 9'h5e == r_count_15_io_out ? io_r_94_b : _GEN_6273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6275 = 9'h5f == r_count_15_io_out ? io_r_95_b : _GEN_6274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6276 = 9'h60 == r_count_15_io_out ? io_r_96_b : _GEN_6275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6277 = 9'h61 == r_count_15_io_out ? io_r_97_b : _GEN_6276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6278 = 9'h62 == r_count_15_io_out ? io_r_98_b : _GEN_6277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6279 = 9'h63 == r_count_15_io_out ? io_r_99_b : _GEN_6278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6280 = 9'h64 == r_count_15_io_out ? io_r_100_b : _GEN_6279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6281 = 9'h65 == r_count_15_io_out ? io_r_101_b : _GEN_6280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6282 = 9'h66 == r_count_15_io_out ? io_r_102_b : _GEN_6281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6283 = 9'h67 == r_count_15_io_out ? io_r_103_b : _GEN_6282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6284 = 9'h68 == r_count_15_io_out ? io_r_104_b : _GEN_6283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6285 = 9'h69 == r_count_15_io_out ? io_r_105_b : _GEN_6284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6286 = 9'h6a == r_count_15_io_out ? io_r_106_b : _GEN_6285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6287 = 9'h6b == r_count_15_io_out ? io_r_107_b : _GEN_6286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6288 = 9'h6c == r_count_15_io_out ? io_r_108_b : _GEN_6287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6289 = 9'h6d == r_count_15_io_out ? io_r_109_b : _GEN_6288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6290 = 9'h6e == r_count_15_io_out ? io_r_110_b : _GEN_6289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6291 = 9'h6f == r_count_15_io_out ? io_r_111_b : _GEN_6290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6292 = 9'h70 == r_count_15_io_out ? io_r_112_b : _GEN_6291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6293 = 9'h71 == r_count_15_io_out ? io_r_113_b : _GEN_6292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6294 = 9'h72 == r_count_15_io_out ? io_r_114_b : _GEN_6293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6295 = 9'h73 == r_count_15_io_out ? io_r_115_b : _GEN_6294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6296 = 9'h74 == r_count_15_io_out ? io_r_116_b : _GEN_6295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6297 = 9'h75 == r_count_15_io_out ? io_r_117_b : _GEN_6296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6298 = 9'h76 == r_count_15_io_out ? io_r_118_b : _GEN_6297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6299 = 9'h77 == r_count_15_io_out ? io_r_119_b : _GEN_6298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6300 = 9'h78 == r_count_15_io_out ? io_r_120_b : _GEN_6299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6301 = 9'h79 == r_count_15_io_out ? io_r_121_b : _GEN_6300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6302 = 9'h7a == r_count_15_io_out ? io_r_122_b : _GEN_6301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6303 = 9'h7b == r_count_15_io_out ? io_r_123_b : _GEN_6302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6304 = 9'h7c == r_count_15_io_out ? io_r_124_b : _GEN_6303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6305 = 9'h7d == r_count_15_io_out ? io_r_125_b : _GEN_6304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6306 = 9'h7e == r_count_15_io_out ? io_r_126_b : _GEN_6305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6307 = 9'h7f == r_count_15_io_out ? io_r_127_b : _GEN_6306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6308 = 9'h80 == r_count_15_io_out ? io_r_128_b : _GEN_6307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6309 = 9'h81 == r_count_15_io_out ? io_r_129_b : _GEN_6308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6310 = 9'h82 == r_count_15_io_out ? io_r_130_b : _GEN_6309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6311 = 9'h83 == r_count_15_io_out ? io_r_131_b : _GEN_6310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6312 = 9'h84 == r_count_15_io_out ? io_r_132_b : _GEN_6311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6313 = 9'h85 == r_count_15_io_out ? io_r_133_b : _GEN_6312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6314 = 9'h86 == r_count_15_io_out ? io_r_134_b : _GEN_6313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6315 = 9'h87 == r_count_15_io_out ? io_r_135_b : _GEN_6314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6316 = 9'h88 == r_count_15_io_out ? io_r_136_b : _GEN_6315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6317 = 9'h89 == r_count_15_io_out ? io_r_137_b : _GEN_6316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6318 = 9'h8a == r_count_15_io_out ? io_r_138_b : _GEN_6317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6319 = 9'h8b == r_count_15_io_out ? io_r_139_b : _GEN_6318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6320 = 9'h8c == r_count_15_io_out ? io_r_140_b : _GEN_6319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6321 = 9'h8d == r_count_15_io_out ? io_r_141_b : _GEN_6320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6322 = 9'h8e == r_count_15_io_out ? io_r_142_b : _GEN_6321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6323 = 9'h8f == r_count_15_io_out ? io_r_143_b : _GEN_6322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6324 = 9'h90 == r_count_15_io_out ? io_r_144_b : _GEN_6323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6325 = 9'h91 == r_count_15_io_out ? io_r_145_b : _GEN_6324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6326 = 9'h92 == r_count_15_io_out ? io_r_146_b : _GEN_6325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6327 = 9'h93 == r_count_15_io_out ? io_r_147_b : _GEN_6326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6328 = 9'h94 == r_count_15_io_out ? io_r_148_b : _GEN_6327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6329 = 9'h95 == r_count_15_io_out ? io_r_149_b : _GEN_6328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6330 = 9'h96 == r_count_15_io_out ? io_r_150_b : _GEN_6329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6331 = 9'h97 == r_count_15_io_out ? io_r_151_b : _GEN_6330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6332 = 9'h98 == r_count_15_io_out ? io_r_152_b : _GEN_6331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6333 = 9'h99 == r_count_15_io_out ? io_r_153_b : _GEN_6332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6334 = 9'h9a == r_count_15_io_out ? io_r_154_b : _GEN_6333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6335 = 9'h9b == r_count_15_io_out ? io_r_155_b : _GEN_6334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6336 = 9'h9c == r_count_15_io_out ? io_r_156_b : _GEN_6335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6337 = 9'h9d == r_count_15_io_out ? io_r_157_b : _GEN_6336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6338 = 9'h9e == r_count_15_io_out ? io_r_158_b : _GEN_6337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6339 = 9'h9f == r_count_15_io_out ? io_r_159_b : _GEN_6338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6340 = 9'ha0 == r_count_15_io_out ? io_r_160_b : _GEN_6339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6341 = 9'ha1 == r_count_15_io_out ? io_r_161_b : _GEN_6340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6342 = 9'ha2 == r_count_15_io_out ? io_r_162_b : _GEN_6341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6343 = 9'ha3 == r_count_15_io_out ? io_r_163_b : _GEN_6342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6344 = 9'ha4 == r_count_15_io_out ? io_r_164_b : _GEN_6343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6345 = 9'ha5 == r_count_15_io_out ? io_r_165_b : _GEN_6344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6346 = 9'ha6 == r_count_15_io_out ? io_r_166_b : _GEN_6345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6347 = 9'ha7 == r_count_15_io_out ? io_r_167_b : _GEN_6346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6348 = 9'ha8 == r_count_15_io_out ? io_r_168_b : _GEN_6347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6349 = 9'ha9 == r_count_15_io_out ? io_r_169_b : _GEN_6348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6350 = 9'haa == r_count_15_io_out ? io_r_170_b : _GEN_6349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6351 = 9'hab == r_count_15_io_out ? io_r_171_b : _GEN_6350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6352 = 9'hac == r_count_15_io_out ? io_r_172_b : _GEN_6351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6353 = 9'had == r_count_15_io_out ? io_r_173_b : _GEN_6352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6354 = 9'hae == r_count_15_io_out ? io_r_174_b : _GEN_6353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6355 = 9'haf == r_count_15_io_out ? io_r_175_b : _GEN_6354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6356 = 9'hb0 == r_count_15_io_out ? io_r_176_b : _GEN_6355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6357 = 9'hb1 == r_count_15_io_out ? io_r_177_b : _GEN_6356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6358 = 9'hb2 == r_count_15_io_out ? io_r_178_b : _GEN_6357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6359 = 9'hb3 == r_count_15_io_out ? io_r_179_b : _GEN_6358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6360 = 9'hb4 == r_count_15_io_out ? io_r_180_b : _GEN_6359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6361 = 9'hb5 == r_count_15_io_out ? io_r_181_b : _GEN_6360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6362 = 9'hb6 == r_count_15_io_out ? io_r_182_b : _GEN_6361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6363 = 9'hb7 == r_count_15_io_out ? io_r_183_b : _GEN_6362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6364 = 9'hb8 == r_count_15_io_out ? io_r_184_b : _GEN_6363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6365 = 9'hb9 == r_count_15_io_out ? io_r_185_b : _GEN_6364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6366 = 9'hba == r_count_15_io_out ? io_r_186_b : _GEN_6365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6367 = 9'hbb == r_count_15_io_out ? io_r_187_b : _GEN_6366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6368 = 9'hbc == r_count_15_io_out ? io_r_188_b : _GEN_6367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6369 = 9'hbd == r_count_15_io_out ? io_r_189_b : _GEN_6368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6370 = 9'hbe == r_count_15_io_out ? io_r_190_b : _GEN_6369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6371 = 9'hbf == r_count_15_io_out ? io_r_191_b : _GEN_6370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6372 = 9'hc0 == r_count_15_io_out ? io_r_192_b : _GEN_6371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6373 = 9'hc1 == r_count_15_io_out ? io_r_193_b : _GEN_6372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6374 = 9'hc2 == r_count_15_io_out ? io_r_194_b : _GEN_6373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6375 = 9'hc3 == r_count_15_io_out ? io_r_195_b : _GEN_6374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6376 = 9'hc4 == r_count_15_io_out ? io_r_196_b : _GEN_6375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6377 = 9'hc5 == r_count_15_io_out ? io_r_197_b : _GEN_6376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6378 = 9'hc6 == r_count_15_io_out ? io_r_198_b : _GEN_6377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6379 = 9'hc7 == r_count_15_io_out ? io_r_199_b : _GEN_6378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6380 = 9'hc8 == r_count_15_io_out ? io_r_200_b : _GEN_6379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6381 = 9'hc9 == r_count_15_io_out ? io_r_201_b : _GEN_6380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6382 = 9'hca == r_count_15_io_out ? io_r_202_b : _GEN_6381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6383 = 9'hcb == r_count_15_io_out ? io_r_203_b : _GEN_6382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6384 = 9'hcc == r_count_15_io_out ? io_r_204_b : _GEN_6383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6385 = 9'hcd == r_count_15_io_out ? io_r_205_b : _GEN_6384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6386 = 9'hce == r_count_15_io_out ? io_r_206_b : _GEN_6385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6387 = 9'hcf == r_count_15_io_out ? io_r_207_b : _GEN_6386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6388 = 9'hd0 == r_count_15_io_out ? io_r_208_b : _GEN_6387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6389 = 9'hd1 == r_count_15_io_out ? io_r_209_b : _GEN_6388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6390 = 9'hd2 == r_count_15_io_out ? io_r_210_b : _GEN_6389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6391 = 9'hd3 == r_count_15_io_out ? io_r_211_b : _GEN_6390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6392 = 9'hd4 == r_count_15_io_out ? io_r_212_b : _GEN_6391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6393 = 9'hd5 == r_count_15_io_out ? io_r_213_b : _GEN_6392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6394 = 9'hd6 == r_count_15_io_out ? io_r_214_b : _GEN_6393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6395 = 9'hd7 == r_count_15_io_out ? io_r_215_b : _GEN_6394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6396 = 9'hd8 == r_count_15_io_out ? io_r_216_b : _GEN_6395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6397 = 9'hd9 == r_count_15_io_out ? io_r_217_b : _GEN_6396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6398 = 9'hda == r_count_15_io_out ? io_r_218_b : _GEN_6397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6399 = 9'hdb == r_count_15_io_out ? io_r_219_b : _GEN_6398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6400 = 9'hdc == r_count_15_io_out ? io_r_220_b : _GEN_6399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6401 = 9'hdd == r_count_15_io_out ? io_r_221_b : _GEN_6400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6402 = 9'hde == r_count_15_io_out ? io_r_222_b : _GEN_6401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6403 = 9'hdf == r_count_15_io_out ? io_r_223_b : _GEN_6402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6404 = 9'he0 == r_count_15_io_out ? io_r_224_b : _GEN_6403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6405 = 9'he1 == r_count_15_io_out ? io_r_225_b : _GEN_6404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6406 = 9'he2 == r_count_15_io_out ? io_r_226_b : _GEN_6405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6407 = 9'he3 == r_count_15_io_out ? io_r_227_b : _GEN_6406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6408 = 9'he4 == r_count_15_io_out ? io_r_228_b : _GEN_6407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6409 = 9'he5 == r_count_15_io_out ? io_r_229_b : _GEN_6408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6410 = 9'he6 == r_count_15_io_out ? io_r_230_b : _GEN_6409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6411 = 9'he7 == r_count_15_io_out ? io_r_231_b : _GEN_6410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6412 = 9'he8 == r_count_15_io_out ? io_r_232_b : _GEN_6411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6413 = 9'he9 == r_count_15_io_out ? io_r_233_b : _GEN_6412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6414 = 9'hea == r_count_15_io_out ? io_r_234_b : _GEN_6413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6415 = 9'heb == r_count_15_io_out ? io_r_235_b : _GEN_6414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6416 = 9'hec == r_count_15_io_out ? io_r_236_b : _GEN_6415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6417 = 9'hed == r_count_15_io_out ? io_r_237_b : _GEN_6416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6418 = 9'hee == r_count_15_io_out ? io_r_238_b : _GEN_6417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6419 = 9'hef == r_count_15_io_out ? io_r_239_b : _GEN_6418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6420 = 9'hf0 == r_count_15_io_out ? io_r_240_b : _GEN_6419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6421 = 9'hf1 == r_count_15_io_out ? io_r_241_b : _GEN_6420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6422 = 9'hf2 == r_count_15_io_out ? io_r_242_b : _GEN_6421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6423 = 9'hf3 == r_count_15_io_out ? io_r_243_b : _GEN_6422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6424 = 9'hf4 == r_count_15_io_out ? io_r_244_b : _GEN_6423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6425 = 9'hf5 == r_count_15_io_out ? io_r_245_b : _GEN_6424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6426 = 9'hf6 == r_count_15_io_out ? io_r_246_b : _GEN_6425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6427 = 9'hf7 == r_count_15_io_out ? io_r_247_b : _GEN_6426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6428 = 9'hf8 == r_count_15_io_out ? io_r_248_b : _GEN_6427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6429 = 9'hf9 == r_count_15_io_out ? io_r_249_b : _GEN_6428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6430 = 9'hfa == r_count_15_io_out ? io_r_250_b : _GEN_6429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6431 = 9'hfb == r_count_15_io_out ? io_r_251_b : _GEN_6430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6432 = 9'hfc == r_count_15_io_out ? io_r_252_b : _GEN_6431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6433 = 9'hfd == r_count_15_io_out ? io_r_253_b : _GEN_6432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6434 = 9'hfe == r_count_15_io_out ? io_r_254_b : _GEN_6433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6435 = 9'hff == r_count_15_io_out ? io_r_255_b : _GEN_6434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6436 = 9'h100 == r_count_15_io_out ? io_r_256_b : _GEN_6435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6437 = 9'h101 == r_count_15_io_out ? io_r_257_b : _GEN_6436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6438 = 9'h102 == r_count_15_io_out ? io_r_258_b : _GEN_6437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6439 = 9'h103 == r_count_15_io_out ? io_r_259_b : _GEN_6438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6440 = 9'h104 == r_count_15_io_out ? io_r_260_b : _GEN_6439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6441 = 9'h105 == r_count_15_io_out ? io_r_261_b : _GEN_6440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6442 = 9'h106 == r_count_15_io_out ? io_r_262_b : _GEN_6441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6443 = 9'h107 == r_count_15_io_out ? io_r_263_b : _GEN_6442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6444 = 9'h108 == r_count_15_io_out ? io_r_264_b : _GEN_6443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6445 = 9'h109 == r_count_15_io_out ? io_r_265_b : _GEN_6444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6446 = 9'h10a == r_count_15_io_out ? io_r_266_b : _GEN_6445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6447 = 9'h10b == r_count_15_io_out ? io_r_267_b : _GEN_6446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6448 = 9'h10c == r_count_15_io_out ? io_r_268_b : _GEN_6447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6449 = 9'h10d == r_count_15_io_out ? io_r_269_b : _GEN_6448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6450 = 9'h10e == r_count_15_io_out ? io_r_270_b : _GEN_6449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6451 = 9'h10f == r_count_15_io_out ? io_r_271_b : _GEN_6450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6452 = 9'h110 == r_count_15_io_out ? io_r_272_b : _GEN_6451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6453 = 9'h111 == r_count_15_io_out ? io_r_273_b : _GEN_6452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6454 = 9'h112 == r_count_15_io_out ? io_r_274_b : _GEN_6453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6455 = 9'h113 == r_count_15_io_out ? io_r_275_b : _GEN_6454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6456 = 9'h114 == r_count_15_io_out ? io_r_276_b : _GEN_6455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6457 = 9'h115 == r_count_15_io_out ? io_r_277_b : _GEN_6456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6458 = 9'h116 == r_count_15_io_out ? io_r_278_b : _GEN_6457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6459 = 9'h117 == r_count_15_io_out ? io_r_279_b : _GEN_6458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6460 = 9'h118 == r_count_15_io_out ? io_r_280_b : _GEN_6459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6461 = 9'h119 == r_count_15_io_out ? io_r_281_b : _GEN_6460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6462 = 9'h11a == r_count_15_io_out ? io_r_282_b : _GEN_6461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6463 = 9'h11b == r_count_15_io_out ? io_r_283_b : _GEN_6462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6464 = 9'h11c == r_count_15_io_out ? io_r_284_b : _GEN_6463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6465 = 9'h11d == r_count_15_io_out ? io_r_285_b : _GEN_6464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6466 = 9'h11e == r_count_15_io_out ? io_r_286_b : _GEN_6465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6467 = 9'h11f == r_count_15_io_out ? io_r_287_b : _GEN_6466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6468 = 9'h120 == r_count_15_io_out ? io_r_288_b : _GEN_6467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6469 = 9'h121 == r_count_15_io_out ? io_r_289_b : _GEN_6468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6470 = 9'h122 == r_count_15_io_out ? io_r_290_b : _GEN_6469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6471 = 9'h123 == r_count_15_io_out ? io_r_291_b : _GEN_6470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6472 = 9'h124 == r_count_15_io_out ? io_r_292_b : _GEN_6471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6473 = 9'h125 == r_count_15_io_out ? io_r_293_b : _GEN_6472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6474 = 9'h126 == r_count_15_io_out ? io_r_294_b : _GEN_6473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6475 = 9'h127 == r_count_15_io_out ? io_r_295_b : _GEN_6474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6476 = 9'h128 == r_count_15_io_out ? io_r_296_b : _GEN_6475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6477 = 9'h129 == r_count_15_io_out ? io_r_297_b : _GEN_6476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6478 = 9'h12a == r_count_15_io_out ? io_r_298_b : _GEN_6477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6479 = 9'h12b == r_count_15_io_out ? io_r_299_b : _GEN_6478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6480 = 9'h12c == r_count_15_io_out ? io_r_300_b : _GEN_6479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6481 = 9'h12d == r_count_15_io_out ? io_r_301_b : _GEN_6480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6482 = 9'h12e == r_count_15_io_out ? io_r_302_b : _GEN_6481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6483 = 9'h12f == r_count_15_io_out ? io_r_303_b : _GEN_6482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6484 = 9'h130 == r_count_15_io_out ? io_r_304_b : _GEN_6483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6485 = 9'h131 == r_count_15_io_out ? io_r_305_b : _GEN_6484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6486 = 9'h132 == r_count_15_io_out ? io_r_306_b : _GEN_6485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6487 = 9'h133 == r_count_15_io_out ? io_r_307_b : _GEN_6486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6488 = 9'h134 == r_count_15_io_out ? io_r_308_b : _GEN_6487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6489 = 9'h135 == r_count_15_io_out ? io_r_309_b : _GEN_6488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6490 = 9'h136 == r_count_15_io_out ? io_r_310_b : _GEN_6489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6491 = 9'h137 == r_count_15_io_out ? io_r_311_b : _GEN_6490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6492 = 9'h138 == r_count_15_io_out ? io_r_312_b : _GEN_6491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6493 = 9'h139 == r_count_15_io_out ? io_r_313_b : _GEN_6492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6494 = 9'h13a == r_count_15_io_out ? io_r_314_b : _GEN_6493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6495 = 9'h13b == r_count_15_io_out ? io_r_315_b : _GEN_6494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6496 = 9'h13c == r_count_15_io_out ? io_r_316_b : _GEN_6495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6497 = 9'h13d == r_count_15_io_out ? io_r_317_b : _GEN_6496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6498 = 9'h13e == r_count_15_io_out ? io_r_318_b : _GEN_6497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6499 = 9'h13f == r_count_15_io_out ? io_r_319_b : _GEN_6498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6500 = 9'h140 == r_count_15_io_out ? io_r_320_b : _GEN_6499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6501 = 9'h141 == r_count_15_io_out ? io_r_321_b : _GEN_6500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6502 = 9'h142 == r_count_15_io_out ? io_r_322_b : _GEN_6501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6503 = 9'h143 == r_count_15_io_out ? io_r_323_b : _GEN_6502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6504 = 9'h144 == r_count_15_io_out ? io_r_324_b : _GEN_6503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6505 = 9'h145 == r_count_15_io_out ? io_r_325_b : _GEN_6504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6506 = 9'h146 == r_count_15_io_out ? io_r_326_b : _GEN_6505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6507 = 9'h147 == r_count_15_io_out ? io_r_327_b : _GEN_6506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6508 = 9'h148 == r_count_15_io_out ? io_r_328_b : _GEN_6507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6509 = 9'h149 == r_count_15_io_out ? io_r_329_b : _GEN_6508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6510 = 9'h14a == r_count_15_io_out ? io_r_330_b : _GEN_6509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6511 = 9'h14b == r_count_15_io_out ? io_r_331_b : _GEN_6510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6512 = 9'h14c == r_count_15_io_out ? io_r_332_b : _GEN_6511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6513 = 9'h14d == r_count_15_io_out ? io_r_333_b : _GEN_6512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6514 = 9'h14e == r_count_15_io_out ? io_r_334_b : _GEN_6513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6515 = 9'h14f == r_count_15_io_out ? io_r_335_b : _GEN_6514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6516 = 9'h150 == r_count_15_io_out ? io_r_336_b : _GEN_6515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6517 = 9'h151 == r_count_15_io_out ? io_r_337_b : _GEN_6516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6518 = 9'h152 == r_count_15_io_out ? io_r_338_b : _GEN_6517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6519 = 9'h153 == r_count_15_io_out ? io_r_339_b : _GEN_6518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6520 = 9'h154 == r_count_15_io_out ? io_r_340_b : _GEN_6519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6521 = 9'h155 == r_count_15_io_out ? io_r_341_b : _GEN_6520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6522 = 9'h156 == r_count_15_io_out ? io_r_342_b : _GEN_6521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6523 = 9'h157 == r_count_15_io_out ? io_r_343_b : _GEN_6522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6524 = 9'h158 == r_count_15_io_out ? io_r_344_b : _GEN_6523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6525 = 9'h159 == r_count_15_io_out ? io_r_345_b : _GEN_6524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6526 = 9'h15a == r_count_15_io_out ? io_r_346_b : _GEN_6525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6527 = 9'h15b == r_count_15_io_out ? io_r_347_b : _GEN_6526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6528 = 9'h15c == r_count_15_io_out ? io_r_348_b : _GEN_6527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6529 = 9'h15d == r_count_15_io_out ? io_r_349_b : _GEN_6528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6530 = 9'h15e == r_count_15_io_out ? io_r_350_b : _GEN_6529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6531 = 9'h15f == r_count_15_io_out ? io_r_351_b : _GEN_6530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6532 = 9'h160 == r_count_15_io_out ? io_r_352_b : _GEN_6531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6533 = 9'h161 == r_count_15_io_out ? io_r_353_b : _GEN_6532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6534 = 9'h162 == r_count_15_io_out ? io_r_354_b : _GEN_6533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6535 = 9'h163 == r_count_15_io_out ? io_r_355_b : _GEN_6534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6536 = 9'h164 == r_count_15_io_out ? io_r_356_b : _GEN_6535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6537 = 9'h165 == r_count_15_io_out ? io_r_357_b : _GEN_6536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6538 = 9'h166 == r_count_15_io_out ? io_r_358_b : _GEN_6537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6539 = 9'h167 == r_count_15_io_out ? io_r_359_b : _GEN_6538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6540 = 9'h168 == r_count_15_io_out ? io_r_360_b : _GEN_6539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6541 = 9'h169 == r_count_15_io_out ? io_r_361_b : _GEN_6540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6542 = 9'h16a == r_count_15_io_out ? io_r_362_b : _GEN_6541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6543 = 9'h16b == r_count_15_io_out ? io_r_363_b : _GEN_6542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6544 = 9'h16c == r_count_15_io_out ? io_r_364_b : _GEN_6543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6545 = 9'h16d == r_count_15_io_out ? io_r_365_b : _GEN_6544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6546 = 9'h16e == r_count_15_io_out ? io_r_366_b : _GEN_6545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6547 = 9'h16f == r_count_15_io_out ? io_r_367_b : _GEN_6546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6548 = 9'h170 == r_count_15_io_out ? io_r_368_b : _GEN_6547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6549 = 9'h171 == r_count_15_io_out ? io_r_369_b : _GEN_6548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6550 = 9'h172 == r_count_15_io_out ? io_r_370_b : _GEN_6549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6551 = 9'h173 == r_count_15_io_out ? io_r_371_b : _GEN_6550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6552 = 9'h174 == r_count_15_io_out ? io_r_372_b : _GEN_6551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6553 = 9'h175 == r_count_15_io_out ? io_r_373_b : _GEN_6552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6554 = 9'h176 == r_count_15_io_out ? io_r_374_b : _GEN_6553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6555 = 9'h177 == r_count_15_io_out ? io_r_375_b : _GEN_6554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6556 = 9'h178 == r_count_15_io_out ? io_r_376_b : _GEN_6555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6557 = 9'h179 == r_count_15_io_out ? io_r_377_b : _GEN_6556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6558 = 9'h17a == r_count_15_io_out ? io_r_378_b : _GEN_6557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6559 = 9'h17b == r_count_15_io_out ? io_r_379_b : _GEN_6558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6560 = 9'h17c == r_count_15_io_out ? io_r_380_b : _GEN_6559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6561 = 9'h17d == r_count_15_io_out ? io_r_381_b : _GEN_6560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6562 = 9'h17e == r_count_15_io_out ? io_r_382_b : _GEN_6561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6563 = 9'h17f == r_count_15_io_out ? io_r_383_b : _GEN_6562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6564 = 9'h180 == r_count_15_io_out ? io_r_384_b : _GEN_6563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6565 = 9'h181 == r_count_15_io_out ? io_r_385_b : _GEN_6564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6566 = 9'h182 == r_count_15_io_out ? io_r_386_b : _GEN_6565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6567 = 9'h183 == r_count_15_io_out ? io_r_387_b : _GEN_6566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6568 = 9'h184 == r_count_15_io_out ? io_r_388_b : _GEN_6567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6569 = 9'h185 == r_count_15_io_out ? io_r_389_b : _GEN_6568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6570 = 9'h186 == r_count_15_io_out ? io_r_390_b : _GEN_6569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6571 = 9'h187 == r_count_15_io_out ? io_r_391_b : _GEN_6570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6572 = 9'h188 == r_count_15_io_out ? io_r_392_b : _GEN_6571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6573 = 9'h189 == r_count_15_io_out ? io_r_393_b : _GEN_6572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6574 = 9'h18a == r_count_15_io_out ? io_r_394_b : _GEN_6573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6575 = 9'h18b == r_count_15_io_out ? io_r_395_b : _GEN_6574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6576 = 9'h18c == r_count_15_io_out ? io_r_396_b : _GEN_6575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6577 = 9'h18d == r_count_15_io_out ? io_r_397_b : _GEN_6576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6578 = 9'h18e == r_count_15_io_out ? io_r_398_b : _GEN_6577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6581 = 9'h1 == r_count_16_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6582 = 9'h2 == r_count_16_io_out ? io_r_2_b : _GEN_6581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6583 = 9'h3 == r_count_16_io_out ? io_r_3_b : _GEN_6582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6584 = 9'h4 == r_count_16_io_out ? io_r_4_b : _GEN_6583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6585 = 9'h5 == r_count_16_io_out ? io_r_5_b : _GEN_6584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6586 = 9'h6 == r_count_16_io_out ? io_r_6_b : _GEN_6585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6587 = 9'h7 == r_count_16_io_out ? io_r_7_b : _GEN_6586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6588 = 9'h8 == r_count_16_io_out ? io_r_8_b : _GEN_6587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6589 = 9'h9 == r_count_16_io_out ? io_r_9_b : _GEN_6588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6590 = 9'ha == r_count_16_io_out ? io_r_10_b : _GEN_6589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6591 = 9'hb == r_count_16_io_out ? io_r_11_b : _GEN_6590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6592 = 9'hc == r_count_16_io_out ? io_r_12_b : _GEN_6591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6593 = 9'hd == r_count_16_io_out ? io_r_13_b : _GEN_6592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6594 = 9'he == r_count_16_io_out ? io_r_14_b : _GEN_6593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6595 = 9'hf == r_count_16_io_out ? io_r_15_b : _GEN_6594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6596 = 9'h10 == r_count_16_io_out ? io_r_16_b : _GEN_6595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6597 = 9'h11 == r_count_16_io_out ? io_r_17_b : _GEN_6596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6598 = 9'h12 == r_count_16_io_out ? io_r_18_b : _GEN_6597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6599 = 9'h13 == r_count_16_io_out ? io_r_19_b : _GEN_6598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6600 = 9'h14 == r_count_16_io_out ? io_r_20_b : _GEN_6599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6601 = 9'h15 == r_count_16_io_out ? io_r_21_b : _GEN_6600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6602 = 9'h16 == r_count_16_io_out ? io_r_22_b : _GEN_6601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6603 = 9'h17 == r_count_16_io_out ? io_r_23_b : _GEN_6602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6604 = 9'h18 == r_count_16_io_out ? io_r_24_b : _GEN_6603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6605 = 9'h19 == r_count_16_io_out ? io_r_25_b : _GEN_6604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6606 = 9'h1a == r_count_16_io_out ? io_r_26_b : _GEN_6605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6607 = 9'h1b == r_count_16_io_out ? io_r_27_b : _GEN_6606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6608 = 9'h1c == r_count_16_io_out ? io_r_28_b : _GEN_6607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6609 = 9'h1d == r_count_16_io_out ? io_r_29_b : _GEN_6608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6610 = 9'h1e == r_count_16_io_out ? io_r_30_b : _GEN_6609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6611 = 9'h1f == r_count_16_io_out ? io_r_31_b : _GEN_6610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6612 = 9'h20 == r_count_16_io_out ? io_r_32_b : _GEN_6611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6613 = 9'h21 == r_count_16_io_out ? io_r_33_b : _GEN_6612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6614 = 9'h22 == r_count_16_io_out ? io_r_34_b : _GEN_6613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6615 = 9'h23 == r_count_16_io_out ? io_r_35_b : _GEN_6614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6616 = 9'h24 == r_count_16_io_out ? io_r_36_b : _GEN_6615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6617 = 9'h25 == r_count_16_io_out ? io_r_37_b : _GEN_6616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6618 = 9'h26 == r_count_16_io_out ? io_r_38_b : _GEN_6617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6619 = 9'h27 == r_count_16_io_out ? io_r_39_b : _GEN_6618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6620 = 9'h28 == r_count_16_io_out ? io_r_40_b : _GEN_6619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6621 = 9'h29 == r_count_16_io_out ? io_r_41_b : _GEN_6620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6622 = 9'h2a == r_count_16_io_out ? io_r_42_b : _GEN_6621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6623 = 9'h2b == r_count_16_io_out ? io_r_43_b : _GEN_6622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6624 = 9'h2c == r_count_16_io_out ? io_r_44_b : _GEN_6623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6625 = 9'h2d == r_count_16_io_out ? io_r_45_b : _GEN_6624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6626 = 9'h2e == r_count_16_io_out ? io_r_46_b : _GEN_6625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6627 = 9'h2f == r_count_16_io_out ? io_r_47_b : _GEN_6626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6628 = 9'h30 == r_count_16_io_out ? io_r_48_b : _GEN_6627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6629 = 9'h31 == r_count_16_io_out ? io_r_49_b : _GEN_6628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6630 = 9'h32 == r_count_16_io_out ? io_r_50_b : _GEN_6629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6631 = 9'h33 == r_count_16_io_out ? io_r_51_b : _GEN_6630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6632 = 9'h34 == r_count_16_io_out ? io_r_52_b : _GEN_6631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6633 = 9'h35 == r_count_16_io_out ? io_r_53_b : _GEN_6632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6634 = 9'h36 == r_count_16_io_out ? io_r_54_b : _GEN_6633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6635 = 9'h37 == r_count_16_io_out ? io_r_55_b : _GEN_6634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6636 = 9'h38 == r_count_16_io_out ? io_r_56_b : _GEN_6635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6637 = 9'h39 == r_count_16_io_out ? io_r_57_b : _GEN_6636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6638 = 9'h3a == r_count_16_io_out ? io_r_58_b : _GEN_6637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6639 = 9'h3b == r_count_16_io_out ? io_r_59_b : _GEN_6638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6640 = 9'h3c == r_count_16_io_out ? io_r_60_b : _GEN_6639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6641 = 9'h3d == r_count_16_io_out ? io_r_61_b : _GEN_6640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6642 = 9'h3e == r_count_16_io_out ? io_r_62_b : _GEN_6641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6643 = 9'h3f == r_count_16_io_out ? io_r_63_b : _GEN_6642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6644 = 9'h40 == r_count_16_io_out ? io_r_64_b : _GEN_6643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6645 = 9'h41 == r_count_16_io_out ? io_r_65_b : _GEN_6644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6646 = 9'h42 == r_count_16_io_out ? io_r_66_b : _GEN_6645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6647 = 9'h43 == r_count_16_io_out ? io_r_67_b : _GEN_6646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6648 = 9'h44 == r_count_16_io_out ? io_r_68_b : _GEN_6647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6649 = 9'h45 == r_count_16_io_out ? io_r_69_b : _GEN_6648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6650 = 9'h46 == r_count_16_io_out ? io_r_70_b : _GEN_6649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6651 = 9'h47 == r_count_16_io_out ? io_r_71_b : _GEN_6650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6652 = 9'h48 == r_count_16_io_out ? io_r_72_b : _GEN_6651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6653 = 9'h49 == r_count_16_io_out ? io_r_73_b : _GEN_6652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6654 = 9'h4a == r_count_16_io_out ? io_r_74_b : _GEN_6653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6655 = 9'h4b == r_count_16_io_out ? io_r_75_b : _GEN_6654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6656 = 9'h4c == r_count_16_io_out ? io_r_76_b : _GEN_6655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6657 = 9'h4d == r_count_16_io_out ? io_r_77_b : _GEN_6656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6658 = 9'h4e == r_count_16_io_out ? io_r_78_b : _GEN_6657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6659 = 9'h4f == r_count_16_io_out ? io_r_79_b : _GEN_6658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6660 = 9'h50 == r_count_16_io_out ? io_r_80_b : _GEN_6659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6661 = 9'h51 == r_count_16_io_out ? io_r_81_b : _GEN_6660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6662 = 9'h52 == r_count_16_io_out ? io_r_82_b : _GEN_6661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6663 = 9'h53 == r_count_16_io_out ? io_r_83_b : _GEN_6662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6664 = 9'h54 == r_count_16_io_out ? io_r_84_b : _GEN_6663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6665 = 9'h55 == r_count_16_io_out ? io_r_85_b : _GEN_6664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6666 = 9'h56 == r_count_16_io_out ? io_r_86_b : _GEN_6665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6667 = 9'h57 == r_count_16_io_out ? io_r_87_b : _GEN_6666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6668 = 9'h58 == r_count_16_io_out ? io_r_88_b : _GEN_6667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6669 = 9'h59 == r_count_16_io_out ? io_r_89_b : _GEN_6668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6670 = 9'h5a == r_count_16_io_out ? io_r_90_b : _GEN_6669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6671 = 9'h5b == r_count_16_io_out ? io_r_91_b : _GEN_6670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6672 = 9'h5c == r_count_16_io_out ? io_r_92_b : _GEN_6671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6673 = 9'h5d == r_count_16_io_out ? io_r_93_b : _GEN_6672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6674 = 9'h5e == r_count_16_io_out ? io_r_94_b : _GEN_6673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6675 = 9'h5f == r_count_16_io_out ? io_r_95_b : _GEN_6674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6676 = 9'h60 == r_count_16_io_out ? io_r_96_b : _GEN_6675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6677 = 9'h61 == r_count_16_io_out ? io_r_97_b : _GEN_6676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6678 = 9'h62 == r_count_16_io_out ? io_r_98_b : _GEN_6677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6679 = 9'h63 == r_count_16_io_out ? io_r_99_b : _GEN_6678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6680 = 9'h64 == r_count_16_io_out ? io_r_100_b : _GEN_6679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6681 = 9'h65 == r_count_16_io_out ? io_r_101_b : _GEN_6680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6682 = 9'h66 == r_count_16_io_out ? io_r_102_b : _GEN_6681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6683 = 9'h67 == r_count_16_io_out ? io_r_103_b : _GEN_6682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6684 = 9'h68 == r_count_16_io_out ? io_r_104_b : _GEN_6683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6685 = 9'h69 == r_count_16_io_out ? io_r_105_b : _GEN_6684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6686 = 9'h6a == r_count_16_io_out ? io_r_106_b : _GEN_6685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6687 = 9'h6b == r_count_16_io_out ? io_r_107_b : _GEN_6686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6688 = 9'h6c == r_count_16_io_out ? io_r_108_b : _GEN_6687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6689 = 9'h6d == r_count_16_io_out ? io_r_109_b : _GEN_6688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6690 = 9'h6e == r_count_16_io_out ? io_r_110_b : _GEN_6689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6691 = 9'h6f == r_count_16_io_out ? io_r_111_b : _GEN_6690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6692 = 9'h70 == r_count_16_io_out ? io_r_112_b : _GEN_6691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6693 = 9'h71 == r_count_16_io_out ? io_r_113_b : _GEN_6692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6694 = 9'h72 == r_count_16_io_out ? io_r_114_b : _GEN_6693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6695 = 9'h73 == r_count_16_io_out ? io_r_115_b : _GEN_6694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6696 = 9'h74 == r_count_16_io_out ? io_r_116_b : _GEN_6695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6697 = 9'h75 == r_count_16_io_out ? io_r_117_b : _GEN_6696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6698 = 9'h76 == r_count_16_io_out ? io_r_118_b : _GEN_6697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6699 = 9'h77 == r_count_16_io_out ? io_r_119_b : _GEN_6698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6700 = 9'h78 == r_count_16_io_out ? io_r_120_b : _GEN_6699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6701 = 9'h79 == r_count_16_io_out ? io_r_121_b : _GEN_6700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6702 = 9'h7a == r_count_16_io_out ? io_r_122_b : _GEN_6701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6703 = 9'h7b == r_count_16_io_out ? io_r_123_b : _GEN_6702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6704 = 9'h7c == r_count_16_io_out ? io_r_124_b : _GEN_6703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6705 = 9'h7d == r_count_16_io_out ? io_r_125_b : _GEN_6704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6706 = 9'h7e == r_count_16_io_out ? io_r_126_b : _GEN_6705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6707 = 9'h7f == r_count_16_io_out ? io_r_127_b : _GEN_6706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6708 = 9'h80 == r_count_16_io_out ? io_r_128_b : _GEN_6707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6709 = 9'h81 == r_count_16_io_out ? io_r_129_b : _GEN_6708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6710 = 9'h82 == r_count_16_io_out ? io_r_130_b : _GEN_6709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6711 = 9'h83 == r_count_16_io_out ? io_r_131_b : _GEN_6710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6712 = 9'h84 == r_count_16_io_out ? io_r_132_b : _GEN_6711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6713 = 9'h85 == r_count_16_io_out ? io_r_133_b : _GEN_6712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6714 = 9'h86 == r_count_16_io_out ? io_r_134_b : _GEN_6713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6715 = 9'h87 == r_count_16_io_out ? io_r_135_b : _GEN_6714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6716 = 9'h88 == r_count_16_io_out ? io_r_136_b : _GEN_6715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6717 = 9'h89 == r_count_16_io_out ? io_r_137_b : _GEN_6716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6718 = 9'h8a == r_count_16_io_out ? io_r_138_b : _GEN_6717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6719 = 9'h8b == r_count_16_io_out ? io_r_139_b : _GEN_6718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6720 = 9'h8c == r_count_16_io_out ? io_r_140_b : _GEN_6719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6721 = 9'h8d == r_count_16_io_out ? io_r_141_b : _GEN_6720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6722 = 9'h8e == r_count_16_io_out ? io_r_142_b : _GEN_6721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6723 = 9'h8f == r_count_16_io_out ? io_r_143_b : _GEN_6722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6724 = 9'h90 == r_count_16_io_out ? io_r_144_b : _GEN_6723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6725 = 9'h91 == r_count_16_io_out ? io_r_145_b : _GEN_6724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6726 = 9'h92 == r_count_16_io_out ? io_r_146_b : _GEN_6725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6727 = 9'h93 == r_count_16_io_out ? io_r_147_b : _GEN_6726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6728 = 9'h94 == r_count_16_io_out ? io_r_148_b : _GEN_6727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6729 = 9'h95 == r_count_16_io_out ? io_r_149_b : _GEN_6728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6730 = 9'h96 == r_count_16_io_out ? io_r_150_b : _GEN_6729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6731 = 9'h97 == r_count_16_io_out ? io_r_151_b : _GEN_6730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6732 = 9'h98 == r_count_16_io_out ? io_r_152_b : _GEN_6731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6733 = 9'h99 == r_count_16_io_out ? io_r_153_b : _GEN_6732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6734 = 9'h9a == r_count_16_io_out ? io_r_154_b : _GEN_6733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6735 = 9'h9b == r_count_16_io_out ? io_r_155_b : _GEN_6734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6736 = 9'h9c == r_count_16_io_out ? io_r_156_b : _GEN_6735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6737 = 9'h9d == r_count_16_io_out ? io_r_157_b : _GEN_6736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6738 = 9'h9e == r_count_16_io_out ? io_r_158_b : _GEN_6737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6739 = 9'h9f == r_count_16_io_out ? io_r_159_b : _GEN_6738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6740 = 9'ha0 == r_count_16_io_out ? io_r_160_b : _GEN_6739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6741 = 9'ha1 == r_count_16_io_out ? io_r_161_b : _GEN_6740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6742 = 9'ha2 == r_count_16_io_out ? io_r_162_b : _GEN_6741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6743 = 9'ha3 == r_count_16_io_out ? io_r_163_b : _GEN_6742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6744 = 9'ha4 == r_count_16_io_out ? io_r_164_b : _GEN_6743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6745 = 9'ha5 == r_count_16_io_out ? io_r_165_b : _GEN_6744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6746 = 9'ha6 == r_count_16_io_out ? io_r_166_b : _GEN_6745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6747 = 9'ha7 == r_count_16_io_out ? io_r_167_b : _GEN_6746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6748 = 9'ha8 == r_count_16_io_out ? io_r_168_b : _GEN_6747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6749 = 9'ha9 == r_count_16_io_out ? io_r_169_b : _GEN_6748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6750 = 9'haa == r_count_16_io_out ? io_r_170_b : _GEN_6749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6751 = 9'hab == r_count_16_io_out ? io_r_171_b : _GEN_6750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6752 = 9'hac == r_count_16_io_out ? io_r_172_b : _GEN_6751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6753 = 9'had == r_count_16_io_out ? io_r_173_b : _GEN_6752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6754 = 9'hae == r_count_16_io_out ? io_r_174_b : _GEN_6753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6755 = 9'haf == r_count_16_io_out ? io_r_175_b : _GEN_6754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6756 = 9'hb0 == r_count_16_io_out ? io_r_176_b : _GEN_6755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6757 = 9'hb1 == r_count_16_io_out ? io_r_177_b : _GEN_6756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6758 = 9'hb2 == r_count_16_io_out ? io_r_178_b : _GEN_6757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6759 = 9'hb3 == r_count_16_io_out ? io_r_179_b : _GEN_6758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6760 = 9'hb4 == r_count_16_io_out ? io_r_180_b : _GEN_6759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6761 = 9'hb5 == r_count_16_io_out ? io_r_181_b : _GEN_6760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6762 = 9'hb6 == r_count_16_io_out ? io_r_182_b : _GEN_6761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6763 = 9'hb7 == r_count_16_io_out ? io_r_183_b : _GEN_6762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6764 = 9'hb8 == r_count_16_io_out ? io_r_184_b : _GEN_6763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6765 = 9'hb9 == r_count_16_io_out ? io_r_185_b : _GEN_6764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6766 = 9'hba == r_count_16_io_out ? io_r_186_b : _GEN_6765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6767 = 9'hbb == r_count_16_io_out ? io_r_187_b : _GEN_6766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6768 = 9'hbc == r_count_16_io_out ? io_r_188_b : _GEN_6767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6769 = 9'hbd == r_count_16_io_out ? io_r_189_b : _GEN_6768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6770 = 9'hbe == r_count_16_io_out ? io_r_190_b : _GEN_6769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6771 = 9'hbf == r_count_16_io_out ? io_r_191_b : _GEN_6770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6772 = 9'hc0 == r_count_16_io_out ? io_r_192_b : _GEN_6771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6773 = 9'hc1 == r_count_16_io_out ? io_r_193_b : _GEN_6772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6774 = 9'hc2 == r_count_16_io_out ? io_r_194_b : _GEN_6773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6775 = 9'hc3 == r_count_16_io_out ? io_r_195_b : _GEN_6774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6776 = 9'hc4 == r_count_16_io_out ? io_r_196_b : _GEN_6775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6777 = 9'hc5 == r_count_16_io_out ? io_r_197_b : _GEN_6776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6778 = 9'hc6 == r_count_16_io_out ? io_r_198_b : _GEN_6777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6779 = 9'hc7 == r_count_16_io_out ? io_r_199_b : _GEN_6778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6780 = 9'hc8 == r_count_16_io_out ? io_r_200_b : _GEN_6779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6781 = 9'hc9 == r_count_16_io_out ? io_r_201_b : _GEN_6780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6782 = 9'hca == r_count_16_io_out ? io_r_202_b : _GEN_6781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6783 = 9'hcb == r_count_16_io_out ? io_r_203_b : _GEN_6782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6784 = 9'hcc == r_count_16_io_out ? io_r_204_b : _GEN_6783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6785 = 9'hcd == r_count_16_io_out ? io_r_205_b : _GEN_6784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6786 = 9'hce == r_count_16_io_out ? io_r_206_b : _GEN_6785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6787 = 9'hcf == r_count_16_io_out ? io_r_207_b : _GEN_6786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6788 = 9'hd0 == r_count_16_io_out ? io_r_208_b : _GEN_6787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6789 = 9'hd1 == r_count_16_io_out ? io_r_209_b : _GEN_6788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6790 = 9'hd2 == r_count_16_io_out ? io_r_210_b : _GEN_6789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6791 = 9'hd3 == r_count_16_io_out ? io_r_211_b : _GEN_6790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6792 = 9'hd4 == r_count_16_io_out ? io_r_212_b : _GEN_6791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6793 = 9'hd5 == r_count_16_io_out ? io_r_213_b : _GEN_6792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6794 = 9'hd6 == r_count_16_io_out ? io_r_214_b : _GEN_6793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6795 = 9'hd7 == r_count_16_io_out ? io_r_215_b : _GEN_6794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6796 = 9'hd8 == r_count_16_io_out ? io_r_216_b : _GEN_6795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6797 = 9'hd9 == r_count_16_io_out ? io_r_217_b : _GEN_6796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6798 = 9'hda == r_count_16_io_out ? io_r_218_b : _GEN_6797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6799 = 9'hdb == r_count_16_io_out ? io_r_219_b : _GEN_6798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6800 = 9'hdc == r_count_16_io_out ? io_r_220_b : _GEN_6799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6801 = 9'hdd == r_count_16_io_out ? io_r_221_b : _GEN_6800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6802 = 9'hde == r_count_16_io_out ? io_r_222_b : _GEN_6801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6803 = 9'hdf == r_count_16_io_out ? io_r_223_b : _GEN_6802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6804 = 9'he0 == r_count_16_io_out ? io_r_224_b : _GEN_6803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6805 = 9'he1 == r_count_16_io_out ? io_r_225_b : _GEN_6804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6806 = 9'he2 == r_count_16_io_out ? io_r_226_b : _GEN_6805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6807 = 9'he3 == r_count_16_io_out ? io_r_227_b : _GEN_6806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6808 = 9'he4 == r_count_16_io_out ? io_r_228_b : _GEN_6807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6809 = 9'he5 == r_count_16_io_out ? io_r_229_b : _GEN_6808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6810 = 9'he6 == r_count_16_io_out ? io_r_230_b : _GEN_6809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6811 = 9'he7 == r_count_16_io_out ? io_r_231_b : _GEN_6810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6812 = 9'he8 == r_count_16_io_out ? io_r_232_b : _GEN_6811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6813 = 9'he9 == r_count_16_io_out ? io_r_233_b : _GEN_6812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6814 = 9'hea == r_count_16_io_out ? io_r_234_b : _GEN_6813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6815 = 9'heb == r_count_16_io_out ? io_r_235_b : _GEN_6814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6816 = 9'hec == r_count_16_io_out ? io_r_236_b : _GEN_6815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6817 = 9'hed == r_count_16_io_out ? io_r_237_b : _GEN_6816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6818 = 9'hee == r_count_16_io_out ? io_r_238_b : _GEN_6817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6819 = 9'hef == r_count_16_io_out ? io_r_239_b : _GEN_6818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6820 = 9'hf0 == r_count_16_io_out ? io_r_240_b : _GEN_6819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6821 = 9'hf1 == r_count_16_io_out ? io_r_241_b : _GEN_6820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6822 = 9'hf2 == r_count_16_io_out ? io_r_242_b : _GEN_6821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6823 = 9'hf3 == r_count_16_io_out ? io_r_243_b : _GEN_6822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6824 = 9'hf4 == r_count_16_io_out ? io_r_244_b : _GEN_6823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6825 = 9'hf5 == r_count_16_io_out ? io_r_245_b : _GEN_6824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6826 = 9'hf6 == r_count_16_io_out ? io_r_246_b : _GEN_6825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6827 = 9'hf7 == r_count_16_io_out ? io_r_247_b : _GEN_6826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6828 = 9'hf8 == r_count_16_io_out ? io_r_248_b : _GEN_6827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6829 = 9'hf9 == r_count_16_io_out ? io_r_249_b : _GEN_6828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6830 = 9'hfa == r_count_16_io_out ? io_r_250_b : _GEN_6829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6831 = 9'hfb == r_count_16_io_out ? io_r_251_b : _GEN_6830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6832 = 9'hfc == r_count_16_io_out ? io_r_252_b : _GEN_6831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6833 = 9'hfd == r_count_16_io_out ? io_r_253_b : _GEN_6832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6834 = 9'hfe == r_count_16_io_out ? io_r_254_b : _GEN_6833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6835 = 9'hff == r_count_16_io_out ? io_r_255_b : _GEN_6834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6836 = 9'h100 == r_count_16_io_out ? io_r_256_b : _GEN_6835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6837 = 9'h101 == r_count_16_io_out ? io_r_257_b : _GEN_6836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6838 = 9'h102 == r_count_16_io_out ? io_r_258_b : _GEN_6837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6839 = 9'h103 == r_count_16_io_out ? io_r_259_b : _GEN_6838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6840 = 9'h104 == r_count_16_io_out ? io_r_260_b : _GEN_6839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6841 = 9'h105 == r_count_16_io_out ? io_r_261_b : _GEN_6840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6842 = 9'h106 == r_count_16_io_out ? io_r_262_b : _GEN_6841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6843 = 9'h107 == r_count_16_io_out ? io_r_263_b : _GEN_6842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6844 = 9'h108 == r_count_16_io_out ? io_r_264_b : _GEN_6843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6845 = 9'h109 == r_count_16_io_out ? io_r_265_b : _GEN_6844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6846 = 9'h10a == r_count_16_io_out ? io_r_266_b : _GEN_6845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6847 = 9'h10b == r_count_16_io_out ? io_r_267_b : _GEN_6846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6848 = 9'h10c == r_count_16_io_out ? io_r_268_b : _GEN_6847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6849 = 9'h10d == r_count_16_io_out ? io_r_269_b : _GEN_6848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6850 = 9'h10e == r_count_16_io_out ? io_r_270_b : _GEN_6849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6851 = 9'h10f == r_count_16_io_out ? io_r_271_b : _GEN_6850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6852 = 9'h110 == r_count_16_io_out ? io_r_272_b : _GEN_6851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6853 = 9'h111 == r_count_16_io_out ? io_r_273_b : _GEN_6852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6854 = 9'h112 == r_count_16_io_out ? io_r_274_b : _GEN_6853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6855 = 9'h113 == r_count_16_io_out ? io_r_275_b : _GEN_6854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6856 = 9'h114 == r_count_16_io_out ? io_r_276_b : _GEN_6855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6857 = 9'h115 == r_count_16_io_out ? io_r_277_b : _GEN_6856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6858 = 9'h116 == r_count_16_io_out ? io_r_278_b : _GEN_6857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6859 = 9'h117 == r_count_16_io_out ? io_r_279_b : _GEN_6858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6860 = 9'h118 == r_count_16_io_out ? io_r_280_b : _GEN_6859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6861 = 9'h119 == r_count_16_io_out ? io_r_281_b : _GEN_6860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6862 = 9'h11a == r_count_16_io_out ? io_r_282_b : _GEN_6861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6863 = 9'h11b == r_count_16_io_out ? io_r_283_b : _GEN_6862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6864 = 9'h11c == r_count_16_io_out ? io_r_284_b : _GEN_6863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6865 = 9'h11d == r_count_16_io_out ? io_r_285_b : _GEN_6864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6866 = 9'h11e == r_count_16_io_out ? io_r_286_b : _GEN_6865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6867 = 9'h11f == r_count_16_io_out ? io_r_287_b : _GEN_6866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6868 = 9'h120 == r_count_16_io_out ? io_r_288_b : _GEN_6867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6869 = 9'h121 == r_count_16_io_out ? io_r_289_b : _GEN_6868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6870 = 9'h122 == r_count_16_io_out ? io_r_290_b : _GEN_6869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6871 = 9'h123 == r_count_16_io_out ? io_r_291_b : _GEN_6870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6872 = 9'h124 == r_count_16_io_out ? io_r_292_b : _GEN_6871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6873 = 9'h125 == r_count_16_io_out ? io_r_293_b : _GEN_6872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6874 = 9'h126 == r_count_16_io_out ? io_r_294_b : _GEN_6873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6875 = 9'h127 == r_count_16_io_out ? io_r_295_b : _GEN_6874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6876 = 9'h128 == r_count_16_io_out ? io_r_296_b : _GEN_6875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6877 = 9'h129 == r_count_16_io_out ? io_r_297_b : _GEN_6876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6878 = 9'h12a == r_count_16_io_out ? io_r_298_b : _GEN_6877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6879 = 9'h12b == r_count_16_io_out ? io_r_299_b : _GEN_6878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6880 = 9'h12c == r_count_16_io_out ? io_r_300_b : _GEN_6879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6881 = 9'h12d == r_count_16_io_out ? io_r_301_b : _GEN_6880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6882 = 9'h12e == r_count_16_io_out ? io_r_302_b : _GEN_6881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6883 = 9'h12f == r_count_16_io_out ? io_r_303_b : _GEN_6882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6884 = 9'h130 == r_count_16_io_out ? io_r_304_b : _GEN_6883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6885 = 9'h131 == r_count_16_io_out ? io_r_305_b : _GEN_6884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6886 = 9'h132 == r_count_16_io_out ? io_r_306_b : _GEN_6885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6887 = 9'h133 == r_count_16_io_out ? io_r_307_b : _GEN_6886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6888 = 9'h134 == r_count_16_io_out ? io_r_308_b : _GEN_6887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6889 = 9'h135 == r_count_16_io_out ? io_r_309_b : _GEN_6888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6890 = 9'h136 == r_count_16_io_out ? io_r_310_b : _GEN_6889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6891 = 9'h137 == r_count_16_io_out ? io_r_311_b : _GEN_6890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6892 = 9'h138 == r_count_16_io_out ? io_r_312_b : _GEN_6891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6893 = 9'h139 == r_count_16_io_out ? io_r_313_b : _GEN_6892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6894 = 9'h13a == r_count_16_io_out ? io_r_314_b : _GEN_6893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6895 = 9'h13b == r_count_16_io_out ? io_r_315_b : _GEN_6894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6896 = 9'h13c == r_count_16_io_out ? io_r_316_b : _GEN_6895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6897 = 9'h13d == r_count_16_io_out ? io_r_317_b : _GEN_6896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6898 = 9'h13e == r_count_16_io_out ? io_r_318_b : _GEN_6897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6899 = 9'h13f == r_count_16_io_out ? io_r_319_b : _GEN_6898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6900 = 9'h140 == r_count_16_io_out ? io_r_320_b : _GEN_6899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6901 = 9'h141 == r_count_16_io_out ? io_r_321_b : _GEN_6900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6902 = 9'h142 == r_count_16_io_out ? io_r_322_b : _GEN_6901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6903 = 9'h143 == r_count_16_io_out ? io_r_323_b : _GEN_6902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6904 = 9'h144 == r_count_16_io_out ? io_r_324_b : _GEN_6903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6905 = 9'h145 == r_count_16_io_out ? io_r_325_b : _GEN_6904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6906 = 9'h146 == r_count_16_io_out ? io_r_326_b : _GEN_6905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6907 = 9'h147 == r_count_16_io_out ? io_r_327_b : _GEN_6906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6908 = 9'h148 == r_count_16_io_out ? io_r_328_b : _GEN_6907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6909 = 9'h149 == r_count_16_io_out ? io_r_329_b : _GEN_6908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6910 = 9'h14a == r_count_16_io_out ? io_r_330_b : _GEN_6909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6911 = 9'h14b == r_count_16_io_out ? io_r_331_b : _GEN_6910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6912 = 9'h14c == r_count_16_io_out ? io_r_332_b : _GEN_6911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6913 = 9'h14d == r_count_16_io_out ? io_r_333_b : _GEN_6912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6914 = 9'h14e == r_count_16_io_out ? io_r_334_b : _GEN_6913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6915 = 9'h14f == r_count_16_io_out ? io_r_335_b : _GEN_6914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6916 = 9'h150 == r_count_16_io_out ? io_r_336_b : _GEN_6915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6917 = 9'h151 == r_count_16_io_out ? io_r_337_b : _GEN_6916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6918 = 9'h152 == r_count_16_io_out ? io_r_338_b : _GEN_6917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6919 = 9'h153 == r_count_16_io_out ? io_r_339_b : _GEN_6918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6920 = 9'h154 == r_count_16_io_out ? io_r_340_b : _GEN_6919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6921 = 9'h155 == r_count_16_io_out ? io_r_341_b : _GEN_6920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6922 = 9'h156 == r_count_16_io_out ? io_r_342_b : _GEN_6921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6923 = 9'h157 == r_count_16_io_out ? io_r_343_b : _GEN_6922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6924 = 9'h158 == r_count_16_io_out ? io_r_344_b : _GEN_6923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6925 = 9'h159 == r_count_16_io_out ? io_r_345_b : _GEN_6924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6926 = 9'h15a == r_count_16_io_out ? io_r_346_b : _GEN_6925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6927 = 9'h15b == r_count_16_io_out ? io_r_347_b : _GEN_6926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6928 = 9'h15c == r_count_16_io_out ? io_r_348_b : _GEN_6927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6929 = 9'h15d == r_count_16_io_out ? io_r_349_b : _GEN_6928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6930 = 9'h15e == r_count_16_io_out ? io_r_350_b : _GEN_6929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6931 = 9'h15f == r_count_16_io_out ? io_r_351_b : _GEN_6930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6932 = 9'h160 == r_count_16_io_out ? io_r_352_b : _GEN_6931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6933 = 9'h161 == r_count_16_io_out ? io_r_353_b : _GEN_6932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6934 = 9'h162 == r_count_16_io_out ? io_r_354_b : _GEN_6933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6935 = 9'h163 == r_count_16_io_out ? io_r_355_b : _GEN_6934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6936 = 9'h164 == r_count_16_io_out ? io_r_356_b : _GEN_6935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6937 = 9'h165 == r_count_16_io_out ? io_r_357_b : _GEN_6936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6938 = 9'h166 == r_count_16_io_out ? io_r_358_b : _GEN_6937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6939 = 9'h167 == r_count_16_io_out ? io_r_359_b : _GEN_6938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6940 = 9'h168 == r_count_16_io_out ? io_r_360_b : _GEN_6939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6941 = 9'h169 == r_count_16_io_out ? io_r_361_b : _GEN_6940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6942 = 9'h16a == r_count_16_io_out ? io_r_362_b : _GEN_6941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6943 = 9'h16b == r_count_16_io_out ? io_r_363_b : _GEN_6942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6944 = 9'h16c == r_count_16_io_out ? io_r_364_b : _GEN_6943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6945 = 9'h16d == r_count_16_io_out ? io_r_365_b : _GEN_6944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6946 = 9'h16e == r_count_16_io_out ? io_r_366_b : _GEN_6945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6947 = 9'h16f == r_count_16_io_out ? io_r_367_b : _GEN_6946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6948 = 9'h170 == r_count_16_io_out ? io_r_368_b : _GEN_6947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6949 = 9'h171 == r_count_16_io_out ? io_r_369_b : _GEN_6948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6950 = 9'h172 == r_count_16_io_out ? io_r_370_b : _GEN_6949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6951 = 9'h173 == r_count_16_io_out ? io_r_371_b : _GEN_6950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6952 = 9'h174 == r_count_16_io_out ? io_r_372_b : _GEN_6951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6953 = 9'h175 == r_count_16_io_out ? io_r_373_b : _GEN_6952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6954 = 9'h176 == r_count_16_io_out ? io_r_374_b : _GEN_6953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6955 = 9'h177 == r_count_16_io_out ? io_r_375_b : _GEN_6954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6956 = 9'h178 == r_count_16_io_out ? io_r_376_b : _GEN_6955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6957 = 9'h179 == r_count_16_io_out ? io_r_377_b : _GEN_6956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6958 = 9'h17a == r_count_16_io_out ? io_r_378_b : _GEN_6957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6959 = 9'h17b == r_count_16_io_out ? io_r_379_b : _GEN_6958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6960 = 9'h17c == r_count_16_io_out ? io_r_380_b : _GEN_6959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6961 = 9'h17d == r_count_16_io_out ? io_r_381_b : _GEN_6960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6962 = 9'h17e == r_count_16_io_out ? io_r_382_b : _GEN_6961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6963 = 9'h17f == r_count_16_io_out ? io_r_383_b : _GEN_6962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6964 = 9'h180 == r_count_16_io_out ? io_r_384_b : _GEN_6963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6965 = 9'h181 == r_count_16_io_out ? io_r_385_b : _GEN_6964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6966 = 9'h182 == r_count_16_io_out ? io_r_386_b : _GEN_6965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6967 = 9'h183 == r_count_16_io_out ? io_r_387_b : _GEN_6966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6968 = 9'h184 == r_count_16_io_out ? io_r_388_b : _GEN_6967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6969 = 9'h185 == r_count_16_io_out ? io_r_389_b : _GEN_6968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6970 = 9'h186 == r_count_16_io_out ? io_r_390_b : _GEN_6969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6971 = 9'h187 == r_count_16_io_out ? io_r_391_b : _GEN_6970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6972 = 9'h188 == r_count_16_io_out ? io_r_392_b : _GEN_6971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6973 = 9'h189 == r_count_16_io_out ? io_r_393_b : _GEN_6972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6974 = 9'h18a == r_count_16_io_out ? io_r_394_b : _GEN_6973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6975 = 9'h18b == r_count_16_io_out ? io_r_395_b : _GEN_6974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6976 = 9'h18c == r_count_16_io_out ? io_r_396_b : _GEN_6975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6977 = 9'h18d == r_count_16_io_out ? io_r_397_b : _GEN_6976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6978 = 9'h18e == r_count_16_io_out ? io_r_398_b : _GEN_6977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6981 = 9'h1 == r_count_17_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6982 = 9'h2 == r_count_17_io_out ? io_r_2_b : _GEN_6981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6983 = 9'h3 == r_count_17_io_out ? io_r_3_b : _GEN_6982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6984 = 9'h4 == r_count_17_io_out ? io_r_4_b : _GEN_6983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6985 = 9'h5 == r_count_17_io_out ? io_r_5_b : _GEN_6984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6986 = 9'h6 == r_count_17_io_out ? io_r_6_b : _GEN_6985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6987 = 9'h7 == r_count_17_io_out ? io_r_7_b : _GEN_6986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6988 = 9'h8 == r_count_17_io_out ? io_r_8_b : _GEN_6987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6989 = 9'h9 == r_count_17_io_out ? io_r_9_b : _GEN_6988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6990 = 9'ha == r_count_17_io_out ? io_r_10_b : _GEN_6989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6991 = 9'hb == r_count_17_io_out ? io_r_11_b : _GEN_6990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6992 = 9'hc == r_count_17_io_out ? io_r_12_b : _GEN_6991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6993 = 9'hd == r_count_17_io_out ? io_r_13_b : _GEN_6992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6994 = 9'he == r_count_17_io_out ? io_r_14_b : _GEN_6993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6995 = 9'hf == r_count_17_io_out ? io_r_15_b : _GEN_6994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6996 = 9'h10 == r_count_17_io_out ? io_r_16_b : _GEN_6995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6997 = 9'h11 == r_count_17_io_out ? io_r_17_b : _GEN_6996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6998 = 9'h12 == r_count_17_io_out ? io_r_18_b : _GEN_6997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6999 = 9'h13 == r_count_17_io_out ? io_r_19_b : _GEN_6998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7000 = 9'h14 == r_count_17_io_out ? io_r_20_b : _GEN_6999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7001 = 9'h15 == r_count_17_io_out ? io_r_21_b : _GEN_7000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7002 = 9'h16 == r_count_17_io_out ? io_r_22_b : _GEN_7001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7003 = 9'h17 == r_count_17_io_out ? io_r_23_b : _GEN_7002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7004 = 9'h18 == r_count_17_io_out ? io_r_24_b : _GEN_7003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7005 = 9'h19 == r_count_17_io_out ? io_r_25_b : _GEN_7004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7006 = 9'h1a == r_count_17_io_out ? io_r_26_b : _GEN_7005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7007 = 9'h1b == r_count_17_io_out ? io_r_27_b : _GEN_7006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7008 = 9'h1c == r_count_17_io_out ? io_r_28_b : _GEN_7007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7009 = 9'h1d == r_count_17_io_out ? io_r_29_b : _GEN_7008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7010 = 9'h1e == r_count_17_io_out ? io_r_30_b : _GEN_7009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7011 = 9'h1f == r_count_17_io_out ? io_r_31_b : _GEN_7010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7012 = 9'h20 == r_count_17_io_out ? io_r_32_b : _GEN_7011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7013 = 9'h21 == r_count_17_io_out ? io_r_33_b : _GEN_7012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7014 = 9'h22 == r_count_17_io_out ? io_r_34_b : _GEN_7013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7015 = 9'h23 == r_count_17_io_out ? io_r_35_b : _GEN_7014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7016 = 9'h24 == r_count_17_io_out ? io_r_36_b : _GEN_7015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7017 = 9'h25 == r_count_17_io_out ? io_r_37_b : _GEN_7016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7018 = 9'h26 == r_count_17_io_out ? io_r_38_b : _GEN_7017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7019 = 9'h27 == r_count_17_io_out ? io_r_39_b : _GEN_7018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7020 = 9'h28 == r_count_17_io_out ? io_r_40_b : _GEN_7019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7021 = 9'h29 == r_count_17_io_out ? io_r_41_b : _GEN_7020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7022 = 9'h2a == r_count_17_io_out ? io_r_42_b : _GEN_7021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7023 = 9'h2b == r_count_17_io_out ? io_r_43_b : _GEN_7022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7024 = 9'h2c == r_count_17_io_out ? io_r_44_b : _GEN_7023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7025 = 9'h2d == r_count_17_io_out ? io_r_45_b : _GEN_7024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7026 = 9'h2e == r_count_17_io_out ? io_r_46_b : _GEN_7025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7027 = 9'h2f == r_count_17_io_out ? io_r_47_b : _GEN_7026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7028 = 9'h30 == r_count_17_io_out ? io_r_48_b : _GEN_7027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7029 = 9'h31 == r_count_17_io_out ? io_r_49_b : _GEN_7028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7030 = 9'h32 == r_count_17_io_out ? io_r_50_b : _GEN_7029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7031 = 9'h33 == r_count_17_io_out ? io_r_51_b : _GEN_7030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7032 = 9'h34 == r_count_17_io_out ? io_r_52_b : _GEN_7031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7033 = 9'h35 == r_count_17_io_out ? io_r_53_b : _GEN_7032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7034 = 9'h36 == r_count_17_io_out ? io_r_54_b : _GEN_7033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7035 = 9'h37 == r_count_17_io_out ? io_r_55_b : _GEN_7034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7036 = 9'h38 == r_count_17_io_out ? io_r_56_b : _GEN_7035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7037 = 9'h39 == r_count_17_io_out ? io_r_57_b : _GEN_7036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7038 = 9'h3a == r_count_17_io_out ? io_r_58_b : _GEN_7037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7039 = 9'h3b == r_count_17_io_out ? io_r_59_b : _GEN_7038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7040 = 9'h3c == r_count_17_io_out ? io_r_60_b : _GEN_7039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7041 = 9'h3d == r_count_17_io_out ? io_r_61_b : _GEN_7040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7042 = 9'h3e == r_count_17_io_out ? io_r_62_b : _GEN_7041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7043 = 9'h3f == r_count_17_io_out ? io_r_63_b : _GEN_7042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7044 = 9'h40 == r_count_17_io_out ? io_r_64_b : _GEN_7043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7045 = 9'h41 == r_count_17_io_out ? io_r_65_b : _GEN_7044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7046 = 9'h42 == r_count_17_io_out ? io_r_66_b : _GEN_7045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7047 = 9'h43 == r_count_17_io_out ? io_r_67_b : _GEN_7046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7048 = 9'h44 == r_count_17_io_out ? io_r_68_b : _GEN_7047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7049 = 9'h45 == r_count_17_io_out ? io_r_69_b : _GEN_7048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7050 = 9'h46 == r_count_17_io_out ? io_r_70_b : _GEN_7049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7051 = 9'h47 == r_count_17_io_out ? io_r_71_b : _GEN_7050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7052 = 9'h48 == r_count_17_io_out ? io_r_72_b : _GEN_7051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7053 = 9'h49 == r_count_17_io_out ? io_r_73_b : _GEN_7052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7054 = 9'h4a == r_count_17_io_out ? io_r_74_b : _GEN_7053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7055 = 9'h4b == r_count_17_io_out ? io_r_75_b : _GEN_7054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7056 = 9'h4c == r_count_17_io_out ? io_r_76_b : _GEN_7055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7057 = 9'h4d == r_count_17_io_out ? io_r_77_b : _GEN_7056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7058 = 9'h4e == r_count_17_io_out ? io_r_78_b : _GEN_7057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7059 = 9'h4f == r_count_17_io_out ? io_r_79_b : _GEN_7058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7060 = 9'h50 == r_count_17_io_out ? io_r_80_b : _GEN_7059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7061 = 9'h51 == r_count_17_io_out ? io_r_81_b : _GEN_7060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7062 = 9'h52 == r_count_17_io_out ? io_r_82_b : _GEN_7061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7063 = 9'h53 == r_count_17_io_out ? io_r_83_b : _GEN_7062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7064 = 9'h54 == r_count_17_io_out ? io_r_84_b : _GEN_7063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7065 = 9'h55 == r_count_17_io_out ? io_r_85_b : _GEN_7064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7066 = 9'h56 == r_count_17_io_out ? io_r_86_b : _GEN_7065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7067 = 9'h57 == r_count_17_io_out ? io_r_87_b : _GEN_7066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7068 = 9'h58 == r_count_17_io_out ? io_r_88_b : _GEN_7067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7069 = 9'h59 == r_count_17_io_out ? io_r_89_b : _GEN_7068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7070 = 9'h5a == r_count_17_io_out ? io_r_90_b : _GEN_7069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7071 = 9'h5b == r_count_17_io_out ? io_r_91_b : _GEN_7070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7072 = 9'h5c == r_count_17_io_out ? io_r_92_b : _GEN_7071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7073 = 9'h5d == r_count_17_io_out ? io_r_93_b : _GEN_7072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7074 = 9'h5e == r_count_17_io_out ? io_r_94_b : _GEN_7073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7075 = 9'h5f == r_count_17_io_out ? io_r_95_b : _GEN_7074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7076 = 9'h60 == r_count_17_io_out ? io_r_96_b : _GEN_7075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7077 = 9'h61 == r_count_17_io_out ? io_r_97_b : _GEN_7076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7078 = 9'h62 == r_count_17_io_out ? io_r_98_b : _GEN_7077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7079 = 9'h63 == r_count_17_io_out ? io_r_99_b : _GEN_7078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7080 = 9'h64 == r_count_17_io_out ? io_r_100_b : _GEN_7079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7081 = 9'h65 == r_count_17_io_out ? io_r_101_b : _GEN_7080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7082 = 9'h66 == r_count_17_io_out ? io_r_102_b : _GEN_7081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7083 = 9'h67 == r_count_17_io_out ? io_r_103_b : _GEN_7082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7084 = 9'h68 == r_count_17_io_out ? io_r_104_b : _GEN_7083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7085 = 9'h69 == r_count_17_io_out ? io_r_105_b : _GEN_7084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7086 = 9'h6a == r_count_17_io_out ? io_r_106_b : _GEN_7085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7087 = 9'h6b == r_count_17_io_out ? io_r_107_b : _GEN_7086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7088 = 9'h6c == r_count_17_io_out ? io_r_108_b : _GEN_7087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7089 = 9'h6d == r_count_17_io_out ? io_r_109_b : _GEN_7088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7090 = 9'h6e == r_count_17_io_out ? io_r_110_b : _GEN_7089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7091 = 9'h6f == r_count_17_io_out ? io_r_111_b : _GEN_7090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7092 = 9'h70 == r_count_17_io_out ? io_r_112_b : _GEN_7091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7093 = 9'h71 == r_count_17_io_out ? io_r_113_b : _GEN_7092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7094 = 9'h72 == r_count_17_io_out ? io_r_114_b : _GEN_7093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7095 = 9'h73 == r_count_17_io_out ? io_r_115_b : _GEN_7094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7096 = 9'h74 == r_count_17_io_out ? io_r_116_b : _GEN_7095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7097 = 9'h75 == r_count_17_io_out ? io_r_117_b : _GEN_7096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7098 = 9'h76 == r_count_17_io_out ? io_r_118_b : _GEN_7097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7099 = 9'h77 == r_count_17_io_out ? io_r_119_b : _GEN_7098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7100 = 9'h78 == r_count_17_io_out ? io_r_120_b : _GEN_7099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7101 = 9'h79 == r_count_17_io_out ? io_r_121_b : _GEN_7100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7102 = 9'h7a == r_count_17_io_out ? io_r_122_b : _GEN_7101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7103 = 9'h7b == r_count_17_io_out ? io_r_123_b : _GEN_7102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7104 = 9'h7c == r_count_17_io_out ? io_r_124_b : _GEN_7103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7105 = 9'h7d == r_count_17_io_out ? io_r_125_b : _GEN_7104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7106 = 9'h7e == r_count_17_io_out ? io_r_126_b : _GEN_7105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7107 = 9'h7f == r_count_17_io_out ? io_r_127_b : _GEN_7106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7108 = 9'h80 == r_count_17_io_out ? io_r_128_b : _GEN_7107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7109 = 9'h81 == r_count_17_io_out ? io_r_129_b : _GEN_7108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7110 = 9'h82 == r_count_17_io_out ? io_r_130_b : _GEN_7109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7111 = 9'h83 == r_count_17_io_out ? io_r_131_b : _GEN_7110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7112 = 9'h84 == r_count_17_io_out ? io_r_132_b : _GEN_7111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7113 = 9'h85 == r_count_17_io_out ? io_r_133_b : _GEN_7112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7114 = 9'h86 == r_count_17_io_out ? io_r_134_b : _GEN_7113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7115 = 9'h87 == r_count_17_io_out ? io_r_135_b : _GEN_7114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7116 = 9'h88 == r_count_17_io_out ? io_r_136_b : _GEN_7115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7117 = 9'h89 == r_count_17_io_out ? io_r_137_b : _GEN_7116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7118 = 9'h8a == r_count_17_io_out ? io_r_138_b : _GEN_7117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7119 = 9'h8b == r_count_17_io_out ? io_r_139_b : _GEN_7118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7120 = 9'h8c == r_count_17_io_out ? io_r_140_b : _GEN_7119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7121 = 9'h8d == r_count_17_io_out ? io_r_141_b : _GEN_7120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7122 = 9'h8e == r_count_17_io_out ? io_r_142_b : _GEN_7121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7123 = 9'h8f == r_count_17_io_out ? io_r_143_b : _GEN_7122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7124 = 9'h90 == r_count_17_io_out ? io_r_144_b : _GEN_7123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7125 = 9'h91 == r_count_17_io_out ? io_r_145_b : _GEN_7124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7126 = 9'h92 == r_count_17_io_out ? io_r_146_b : _GEN_7125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7127 = 9'h93 == r_count_17_io_out ? io_r_147_b : _GEN_7126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7128 = 9'h94 == r_count_17_io_out ? io_r_148_b : _GEN_7127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7129 = 9'h95 == r_count_17_io_out ? io_r_149_b : _GEN_7128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7130 = 9'h96 == r_count_17_io_out ? io_r_150_b : _GEN_7129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7131 = 9'h97 == r_count_17_io_out ? io_r_151_b : _GEN_7130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7132 = 9'h98 == r_count_17_io_out ? io_r_152_b : _GEN_7131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7133 = 9'h99 == r_count_17_io_out ? io_r_153_b : _GEN_7132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7134 = 9'h9a == r_count_17_io_out ? io_r_154_b : _GEN_7133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7135 = 9'h9b == r_count_17_io_out ? io_r_155_b : _GEN_7134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7136 = 9'h9c == r_count_17_io_out ? io_r_156_b : _GEN_7135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7137 = 9'h9d == r_count_17_io_out ? io_r_157_b : _GEN_7136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7138 = 9'h9e == r_count_17_io_out ? io_r_158_b : _GEN_7137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7139 = 9'h9f == r_count_17_io_out ? io_r_159_b : _GEN_7138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7140 = 9'ha0 == r_count_17_io_out ? io_r_160_b : _GEN_7139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7141 = 9'ha1 == r_count_17_io_out ? io_r_161_b : _GEN_7140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7142 = 9'ha2 == r_count_17_io_out ? io_r_162_b : _GEN_7141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7143 = 9'ha3 == r_count_17_io_out ? io_r_163_b : _GEN_7142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7144 = 9'ha4 == r_count_17_io_out ? io_r_164_b : _GEN_7143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7145 = 9'ha5 == r_count_17_io_out ? io_r_165_b : _GEN_7144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7146 = 9'ha6 == r_count_17_io_out ? io_r_166_b : _GEN_7145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7147 = 9'ha7 == r_count_17_io_out ? io_r_167_b : _GEN_7146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7148 = 9'ha8 == r_count_17_io_out ? io_r_168_b : _GEN_7147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7149 = 9'ha9 == r_count_17_io_out ? io_r_169_b : _GEN_7148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7150 = 9'haa == r_count_17_io_out ? io_r_170_b : _GEN_7149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7151 = 9'hab == r_count_17_io_out ? io_r_171_b : _GEN_7150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7152 = 9'hac == r_count_17_io_out ? io_r_172_b : _GEN_7151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7153 = 9'had == r_count_17_io_out ? io_r_173_b : _GEN_7152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7154 = 9'hae == r_count_17_io_out ? io_r_174_b : _GEN_7153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7155 = 9'haf == r_count_17_io_out ? io_r_175_b : _GEN_7154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7156 = 9'hb0 == r_count_17_io_out ? io_r_176_b : _GEN_7155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7157 = 9'hb1 == r_count_17_io_out ? io_r_177_b : _GEN_7156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7158 = 9'hb2 == r_count_17_io_out ? io_r_178_b : _GEN_7157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7159 = 9'hb3 == r_count_17_io_out ? io_r_179_b : _GEN_7158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7160 = 9'hb4 == r_count_17_io_out ? io_r_180_b : _GEN_7159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7161 = 9'hb5 == r_count_17_io_out ? io_r_181_b : _GEN_7160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7162 = 9'hb6 == r_count_17_io_out ? io_r_182_b : _GEN_7161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7163 = 9'hb7 == r_count_17_io_out ? io_r_183_b : _GEN_7162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7164 = 9'hb8 == r_count_17_io_out ? io_r_184_b : _GEN_7163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7165 = 9'hb9 == r_count_17_io_out ? io_r_185_b : _GEN_7164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7166 = 9'hba == r_count_17_io_out ? io_r_186_b : _GEN_7165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7167 = 9'hbb == r_count_17_io_out ? io_r_187_b : _GEN_7166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7168 = 9'hbc == r_count_17_io_out ? io_r_188_b : _GEN_7167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7169 = 9'hbd == r_count_17_io_out ? io_r_189_b : _GEN_7168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7170 = 9'hbe == r_count_17_io_out ? io_r_190_b : _GEN_7169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7171 = 9'hbf == r_count_17_io_out ? io_r_191_b : _GEN_7170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7172 = 9'hc0 == r_count_17_io_out ? io_r_192_b : _GEN_7171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7173 = 9'hc1 == r_count_17_io_out ? io_r_193_b : _GEN_7172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7174 = 9'hc2 == r_count_17_io_out ? io_r_194_b : _GEN_7173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7175 = 9'hc3 == r_count_17_io_out ? io_r_195_b : _GEN_7174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7176 = 9'hc4 == r_count_17_io_out ? io_r_196_b : _GEN_7175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7177 = 9'hc5 == r_count_17_io_out ? io_r_197_b : _GEN_7176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7178 = 9'hc6 == r_count_17_io_out ? io_r_198_b : _GEN_7177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7179 = 9'hc7 == r_count_17_io_out ? io_r_199_b : _GEN_7178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7180 = 9'hc8 == r_count_17_io_out ? io_r_200_b : _GEN_7179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7181 = 9'hc9 == r_count_17_io_out ? io_r_201_b : _GEN_7180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7182 = 9'hca == r_count_17_io_out ? io_r_202_b : _GEN_7181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7183 = 9'hcb == r_count_17_io_out ? io_r_203_b : _GEN_7182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7184 = 9'hcc == r_count_17_io_out ? io_r_204_b : _GEN_7183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7185 = 9'hcd == r_count_17_io_out ? io_r_205_b : _GEN_7184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7186 = 9'hce == r_count_17_io_out ? io_r_206_b : _GEN_7185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7187 = 9'hcf == r_count_17_io_out ? io_r_207_b : _GEN_7186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7188 = 9'hd0 == r_count_17_io_out ? io_r_208_b : _GEN_7187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7189 = 9'hd1 == r_count_17_io_out ? io_r_209_b : _GEN_7188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7190 = 9'hd2 == r_count_17_io_out ? io_r_210_b : _GEN_7189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7191 = 9'hd3 == r_count_17_io_out ? io_r_211_b : _GEN_7190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7192 = 9'hd4 == r_count_17_io_out ? io_r_212_b : _GEN_7191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7193 = 9'hd5 == r_count_17_io_out ? io_r_213_b : _GEN_7192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7194 = 9'hd6 == r_count_17_io_out ? io_r_214_b : _GEN_7193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7195 = 9'hd7 == r_count_17_io_out ? io_r_215_b : _GEN_7194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7196 = 9'hd8 == r_count_17_io_out ? io_r_216_b : _GEN_7195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7197 = 9'hd9 == r_count_17_io_out ? io_r_217_b : _GEN_7196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7198 = 9'hda == r_count_17_io_out ? io_r_218_b : _GEN_7197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7199 = 9'hdb == r_count_17_io_out ? io_r_219_b : _GEN_7198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7200 = 9'hdc == r_count_17_io_out ? io_r_220_b : _GEN_7199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7201 = 9'hdd == r_count_17_io_out ? io_r_221_b : _GEN_7200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7202 = 9'hde == r_count_17_io_out ? io_r_222_b : _GEN_7201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7203 = 9'hdf == r_count_17_io_out ? io_r_223_b : _GEN_7202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7204 = 9'he0 == r_count_17_io_out ? io_r_224_b : _GEN_7203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7205 = 9'he1 == r_count_17_io_out ? io_r_225_b : _GEN_7204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7206 = 9'he2 == r_count_17_io_out ? io_r_226_b : _GEN_7205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7207 = 9'he3 == r_count_17_io_out ? io_r_227_b : _GEN_7206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7208 = 9'he4 == r_count_17_io_out ? io_r_228_b : _GEN_7207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7209 = 9'he5 == r_count_17_io_out ? io_r_229_b : _GEN_7208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7210 = 9'he6 == r_count_17_io_out ? io_r_230_b : _GEN_7209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7211 = 9'he7 == r_count_17_io_out ? io_r_231_b : _GEN_7210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7212 = 9'he8 == r_count_17_io_out ? io_r_232_b : _GEN_7211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7213 = 9'he9 == r_count_17_io_out ? io_r_233_b : _GEN_7212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7214 = 9'hea == r_count_17_io_out ? io_r_234_b : _GEN_7213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7215 = 9'heb == r_count_17_io_out ? io_r_235_b : _GEN_7214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7216 = 9'hec == r_count_17_io_out ? io_r_236_b : _GEN_7215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7217 = 9'hed == r_count_17_io_out ? io_r_237_b : _GEN_7216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7218 = 9'hee == r_count_17_io_out ? io_r_238_b : _GEN_7217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7219 = 9'hef == r_count_17_io_out ? io_r_239_b : _GEN_7218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7220 = 9'hf0 == r_count_17_io_out ? io_r_240_b : _GEN_7219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7221 = 9'hf1 == r_count_17_io_out ? io_r_241_b : _GEN_7220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7222 = 9'hf2 == r_count_17_io_out ? io_r_242_b : _GEN_7221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7223 = 9'hf3 == r_count_17_io_out ? io_r_243_b : _GEN_7222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7224 = 9'hf4 == r_count_17_io_out ? io_r_244_b : _GEN_7223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7225 = 9'hf5 == r_count_17_io_out ? io_r_245_b : _GEN_7224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7226 = 9'hf6 == r_count_17_io_out ? io_r_246_b : _GEN_7225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7227 = 9'hf7 == r_count_17_io_out ? io_r_247_b : _GEN_7226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7228 = 9'hf8 == r_count_17_io_out ? io_r_248_b : _GEN_7227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7229 = 9'hf9 == r_count_17_io_out ? io_r_249_b : _GEN_7228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7230 = 9'hfa == r_count_17_io_out ? io_r_250_b : _GEN_7229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7231 = 9'hfb == r_count_17_io_out ? io_r_251_b : _GEN_7230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7232 = 9'hfc == r_count_17_io_out ? io_r_252_b : _GEN_7231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7233 = 9'hfd == r_count_17_io_out ? io_r_253_b : _GEN_7232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7234 = 9'hfe == r_count_17_io_out ? io_r_254_b : _GEN_7233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7235 = 9'hff == r_count_17_io_out ? io_r_255_b : _GEN_7234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7236 = 9'h100 == r_count_17_io_out ? io_r_256_b : _GEN_7235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7237 = 9'h101 == r_count_17_io_out ? io_r_257_b : _GEN_7236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7238 = 9'h102 == r_count_17_io_out ? io_r_258_b : _GEN_7237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7239 = 9'h103 == r_count_17_io_out ? io_r_259_b : _GEN_7238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7240 = 9'h104 == r_count_17_io_out ? io_r_260_b : _GEN_7239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7241 = 9'h105 == r_count_17_io_out ? io_r_261_b : _GEN_7240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7242 = 9'h106 == r_count_17_io_out ? io_r_262_b : _GEN_7241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7243 = 9'h107 == r_count_17_io_out ? io_r_263_b : _GEN_7242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7244 = 9'h108 == r_count_17_io_out ? io_r_264_b : _GEN_7243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7245 = 9'h109 == r_count_17_io_out ? io_r_265_b : _GEN_7244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7246 = 9'h10a == r_count_17_io_out ? io_r_266_b : _GEN_7245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7247 = 9'h10b == r_count_17_io_out ? io_r_267_b : _GEN_7246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7248 = 9'h10c == r_count_17_io_out ? io_r_268_b : _GEN_7247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7249 = 9'h10d == r_count_17_io_out ? io_r_269_b : _GEN_7248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7250 = 9'h10e == r_count_17_io_out ? io_r_270_b : _GEN_7249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7251 = 9'h10f == r_count_17_io_out ? io_r_271_b : _GEN_7250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7252 = 9'h110 == r_count_17_io_out ? io_r_272_b : _GEN_7251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7253 = 9'h111 == r_count_17_io_out ? io_r_273_b : _GEN_7252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7254 = 9'h112 == r_count_17_io_out ? io_r_274_b : _GEN_7253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7255 = 9'h113 == r_count_17_io_out ? io_r_275_b : _GEN_7254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7256 = 9'h114 == r_count_17_io_out ? io_r_276_b : _GEN_7255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7257 = 9'h115 == r_count_17_io_out ? io_r_277_b : _GEN_7256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7258 = 9'h116 == r_count_17_io_out ? io_r_278_b : _GEN_7257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7259 = 9'h117 == r_count_17_io_out ? io_r_279_b : _GEN_7258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7260 = 9'h118 == r_count_17_io_out ? io_r_280_b : _GEN_7259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7261 = 9'h119 == r_count_17_io_out ? io_r_281_b : _GEN_7260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7262 = 9'h11a == r_count_17_io_out ? io_r_282_b : _GEN_7261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7263 = 9'h11b == r_count_17_io_out ? io_r_283_b : _GEN_7262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7264 = 9'h11c == r_count_17_io_out ? io_r_284_b : _GEN_7263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7265 = 9'h11d == r_count_17_io_out ? io_r_285_b : _GEN_7264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7266 = 9'h11e == r_count_17_io_out ? io_r_286_b : _GEN_7265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7267 = 9'h11f == r_count_17_io_out ? io_r_287_b : _GEN_7266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7268 = 9'h120 == r_count_17_io_out ? io_r_288_b : _GEN_7267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7269 = 9'h121 == r_count_17_io_out ? io_r_289_b : _GEN_7268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7270 = 9'h122 == r_count_17_io_out ? io_r_290_b : _GEN_7269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7271 = 9'h123 == r_count_17_io_out ? io_r_291_b : _GEN_7270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7272 = 9'h124 == r_count_17_io_out ? io_r_292_b : _GEN_7271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7273 = 9'h125 == r_count_17_io_out ? io_r_293_b : _GEN_7272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7274 = 9'h126 == r_count_17_io_out ? io_r_294_b : _GEN_7273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7275 = 9'h127 == r_count_17_io_out ? io_r_295_b : _GEN_7274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7276 = 9'h128 == r_count_17_io_out ? io_r_296_b : _GEN_7275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7277 = 9'h129 == r_count_17_io_out ? io_r_297_b : _GEN_7276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7278 = 9'h12a == r_count_17_io_out ? io_r_298_b : _GEN_7277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7279 = 9'h12b == r_count_17_io_out ? io_r_299_b : _GEN_7278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7280 = 9'h12c == r_count_17_io_out ? io_r_300_b : _GEN_7279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7281 = 9'h12d == r_count_17_io_out ? io_r_301_b : _GEN_7280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7282 = 9'h12e == r_count_17_io_out ? io_r_302_b : _GEN_7281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7283 = 9'h12f == r_count_17_io_out ? io_r_303_b : _GEN_7282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7284 = 9'h130 == r_count_17_io_out ? io_r_304_b : _GEN_7283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7285 = 9'h131 == r_count_17_io_out ? io_r_305_b : _GEN_7284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7286 = 9'h132 == r_count_17_io_out ? io_r_306_b : _GEN_7285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7287 = 9'h133 == r_count_17_io_out ? io_r_307_b : _GEN_7286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7288 = 9'h134 == r_count_17_io_out ? io_r_308_b : _GEN_7287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7289 = 9'h135 == r_count_17_io_out ? io_r_309_b : _GEN_7288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7290 = 9'h136 == r_count_17_io_out ? io_r_310_b : _GEN_7289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7291 = 9'h137 == r_count_17_io_out ? io_r_311_b : _GEN_7290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7292 = 9'h138 == r_count_17_io_out ? io_r_312_b : _GEN_7291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7293 = 9'h139 == r_count_17_io_out ? io_r_313_b : _GEN_7292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7294 = 9'h13a == r_count_17_io_out ? io_r_314_b : _GEN_7293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7295 = 9'h13b == r_count_17_io_out ? io_r_315_b : _GEN_7294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7296 = 9'h13c == r_count_17_io_out ? io_r_316_b : _GEN_7295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7297 = 9'h13d == r_count_17_io_out ? io_r_317_b : _GEN_7296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7298 = 9'h13e == r_count_17_io_out ? io_r_318_b : _GEN_7297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7299 = 9'h13f == r_count_17_io_out ? io_r_319_b : _GEN_7298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7300 = 9'h140 == r_count_17_io_out ? io_r_320_b : _GEN_7299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7301 = 9'h141 == r_count_17_io_out ? io_r_321_b : _GEN_7300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7302 = 9'h142 == r_count_17_io_out ? io_r_322_b : _GEN_7301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7303 = 9'h143 == r_count_17_io_out ? io_r_323_b : _GEN_7302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7304 = 9'h144 == r_count_17_io_out ? io_r_324_b : _GEN_7303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7305 = 9'h145 == r_count_17_io_out ? io_r_325_b : _GEN_7304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7306 = 9'h146 == r_count_17_io_out ? io_r_326_b : _GEN_7305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7307 = 9'h147 == r_count_17_io_out ? io_r_327_b : _GEN_7306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7308 = 9'h148 == r_count_17_io_out ? io_r_328_b : _GEN_7307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7309 = 9'h149 == r_count_17_io_out ? io_r_329_b : _GEN_7308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7310 = 9'h14a == r_count_17_io_out ? io_r_330_b : _GEN_7309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7311 = 9'h14b == r_count_17_io_out ? io_r_331_b : _GEN_7310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7312 = 9'h14c == r_count_17_io_out ? io_r_332_b : _GEN_7311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7313 = 9'h14d == r_count_17_io_out ? io_r_333_b : _GEN_7312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7314 = 9'h14e == r_count_17_io_out ? io_r_334_b : _GEN_7313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7315 = 9'h14f == r_count_17_io_out ? io_r_335_b : _GEN_7314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7316 = 9'h150 == r_count_17_io_out ? io_r_336_b : _GEN_7315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7317 = 9'h151 == r_count_17_io_out ? io_r_337_b : _GEN_7316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7318 = 9'h152 == r_count_17_io_out ? io_r_338_b : _GEN_7317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7319 = 9'h153 == r_count_17_io_out ? io_r_339_b : _GEN_7318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7320 = 9'h154 == r_count_17_io_out ? io_r_340_b : _GEN_7319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7321 = 9'h155 == r_count_17_io_out ? io_r_341_b : _GEN_7320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7322 = 9'h156 == r_count_17_io_out ? io_r_342_b : _GEN_7321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7323 = 9'h157 == r_count_17_io_out ? io_r_343_b : _GEN_7322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7324 = 9'h158 == r_count_17_io_out ? io_r_344_b : _GEN_7323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7325 = 9'h159 == r_count_17_io_out ? io_r_345_b : _GEN_7324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7326 = 9'h15a == r_count_17_io_out ? io_r_346_b : _GEN_7325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7327 = 9'h15b == r_count_17_io_out ? io_r_347_b : _GEN_7326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7328 = 9'h15c == r_count_17_io_out ? io_r_348_b : _GEN_7327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7329 = 9'h15d == r_count_17_io_out ? io_r_349_b : _GEN_7328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7330 = 9'h15e == r_count_17_io_out ? io_r_350_b : _GEN_7329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7331 = 9'h15f == r_count_17_io_out ? io_r_351_b : _GEN_7330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7332 = 9'h160 == r_count_17_io_out ? io_r_352_b : _GEN_7331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7333 = 9'h161 == r_count_17_io_out ? io_r_353_b : _GEN_7332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7334 = 9'h162 == r_count_17_io_out ? io_r_354_b : _GEN_7333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7335 = 9'h163 == r_count_17_io_out ? io_r_355_b : _GEN_7334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7336 = 9'h164 == r_count_17_io_out ? io_r_356_b : _GEN_7335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7337 = 9'h165 == r_count_17_io_out ? io_r_357_b : _GEN_7336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7338 = 9'h166 == r_count_17_io_out ? io_r_358_b : _GEN_7337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7339 = 9'h167 == r_count_17_io_out ? io_r_359_b : _GEN_7338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7340 = 9'h168 == r_count_17_io_out ? io_r_360_b : _GEN_7339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7341 = 9'h169 == r_count_17_io_out ? io_r_361_b : _GEN_7340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7342 = 9'h16a == r_count_17_io_out ? io_r_362_b : _GEN_7341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7343 = 9'h16b == r_count_17_io_out ? io_r_363_b : _GEN_7342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7344 = 9'h16c == r_count_17_io_out ? io_r_364_b : _GEN_7343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7345 = 9'h16d == r_count_17_io_out ? io_r_365_b : _GEN_7344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7346 = 9'h16e == r_count_17_io_out ? io_r_366_b : _GEN_7345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7347 = 9'h16f == r_count_17_io_out ? io_r_367_b : _GEN_7346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7348 = 9'h170 == r_count_17_io_out ? io_r_368_b : _GEN_7347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7349 = 9'h171 == r_count_17_io_out ? io_r_369_b : _GEN_7348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7350 = 9'h172 == r_count_17_io_out ? io_r_370_b : _GEN_7349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7351 = 9'h173 == r_count_17_io_out ? io_r_371_b : _GEN_7350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7352 = 9'h174 == r_count_17_io_out ? io_r_372_b : _GEN_7351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7353 = 9'h175 == r_count_17_io_out ? io_r_373_b : _GEN_7352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7354 = 9'h176 == r_count_17_io_out ? io_r_374_b : _GEN_7353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7355 = 9'h177 == r_count_17_io_out ? io_r_375_b : _GEN_7354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7356 = 9'h178 == r_count_17_io_out ? io_r_376_b : _GEN_7355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7357 = 9'h179 == r_count_17_io_out ? io_r_377_b : _GEN_7356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7358 = 9'h17a == r_count_17_io_out ? io_r_378_b : _GEN_7357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7359 = 9'h17b == r_count_17_io_out ? io_r_379_b : _GEN_7358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7360 = 9'h17c == r_count_17_io_out ? io_r_380_b : _GEN_7359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7361 = 9'h17d == r_count_17_io_out ? io_r_381_b : _GEN_7360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7362 = 9'h17e == r_count_17_io_out ? io_r_382_b : _GEN_7361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7363 = 9'h17f == r_count_17_io_out ? io_r_383_b : _GEN_7362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7364 = 9'h180 == r_count_17_io_out ? io_r_384_b : _GEN_7363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7365 = 9'h181 == r_count_17_io_out ? io_r_385_b : _GEN_7364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7366 = 9'h182 == r_count_17_io_out ? io_r_386_b : _GEN_7365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7367 = 9'h183 == r_count_17_io_out ? io_r_387_b : _GEN_7366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7368 = 9'h184 == r_count_17_io_out ? io_r_388_b : _GEN_7367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7369 = 9'h185 == r_count_17_io_out ? io_r_389_b : _GEN_7368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7370 = 9'h186 == r_count_17_io_out ? io_r_390_b : _GEN_7369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7371 = 9'h187 == r_count_17_io_out ? io_r_391_b : _GEN_7370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7372 = 9'h188 == r_count_17_io_out ? io_r_392_b : _GEN_7371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7373 = 9'h189 == r_count_17_io_out ? io_r_393_b : _GEN_7372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7374 = 9'h18a == r_count_17_io_out ? io_r_394_b : _GEN_7373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7375 = 9'h18b == r_count_17_io_out ? io_r_395_b : _GEN_7374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7376 = 9'h18c == r_count_17_io_out ? io_r_396_b : _GEN_7375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7377 = 9'h18d == r_count_17_io_out ? io_r_397_b : _GEN_7376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7378 = 9'h18e == r_count_17_io_out ? io_r_398_b : _GEN_7377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7381 = 9'h1 == r_count_18_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7382 = 9'h2 == r_count_18_io_out ? io_r_2_b : _GEN_7381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7383 = 9'h3 == r_count_18_io_out ? io_r_3_b : _GEN_7382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7384 = 9'h4 == r_count_18_io_out ? io_r_4_b : _GEN_7383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7385 = 9'h5 == r_count_18_io_out ? io_r_5_b : _GEN_7384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7386 = 9'h6 == r_count_18_io_out ? io_r_6_b : _GEN_7385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7387 = 9'h7 == r_count_18_io_out ? io_r_7_b : _GEN_7386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7388 = 9'h8 == r_count_18_io_out ? io_r_8_b : _GEN_7387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7389 = 9'h9 == r_count_18_io_out ? io_r_9_b : _GEN_7388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7390 = 9'ha == r_count_18_io_out ? io_r_10_b : _GEN_7389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7391 = 9'hb == r_count_18_io_out ? io_r_11_b : _GEN_7390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7392 = 9'hc == r_count_18_io_out ? io_r_12_b : _GEN_7391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7393 = 9'hd == r_count_18_io_out ? io_r_13_b : _GEN_7392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7394 = 9'he == r_count_18_io_out ? io_r_14_b : _GEN_7393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7395 = 9'hf == r_count_18_io_out ? io_r_15_b : _GEN_7394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7396 = 9'h10 == r_count_18_io_out ? io_r_16_b : _GEN_7395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7397 = 9'h11 == r_count_18_io_out ? io_r_17_b : _GEN_7396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7398 = 9'h12 == r_count_18_io_out ? io_r_18_b : _GEN_7397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7399 = 9'h13 == r_count_18_io_out ? io_r_19_b : _GEN_7398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7400 = 9'h14 == r_count_18_io_out ? io_r_20_b : _GEN_7399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7401 = 9'h15 == r_count_18_io_out ? io_r_21_b : _GEN_7400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7402 = 9'h16 == r_count_18_io_out ? io_r_22_b : _GEN_7401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7403 = 9'h17 == r_count_18_io_out ? io_r_23_b : _GEN_7402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7404 = 9'h18 == r_count_18_io_out ? io_r_24_b : _GEN_7403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7405 = 9'h19 == r_count_18_io_out ? io_r_25_b : _GEN_7404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7406 = 9'h1a == r_count_18_io_out ? io_r_26_b : _GEN_7405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7407 = 9'h1b == r_count_18_io_out ? io_r_27_b : _GEN_7406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7408 = 9'h1c == r_count_18_io_out ? io_r_28_b : _GEN_7407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7409 = 9'h1d == r_count_18_io_out ? io_r_29_b : _GEN_7408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7410 = 9'h1e == r_count_18_io_out ? io_r_30_b : _GEN_7409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7411 = 9'h1f == r_count_18_io_out ? io_r_31_b : _GEN_7410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7412 = 9'h20 == r_count_18_io_out ? io_r_32_b : _GEN_7411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7413 = 9'h21 == r_count_18_io_out ? io_r_33_b : _GEN_7412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7414 = 9'h22 == r_count_18_io_out ? io_r_34_b : _GEN_7413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7415 = 9'h23 == r_count_18_io_out ? io_r_35_b : _GEN_7414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7416 = 9'h24 == r_count_18_io_out ? io_r_36_b : _GEN_7415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7417 = 9'h25 == r_count_18_io_out ? io_r_37_b : _GEN_7416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7418 = 9'h26 == r_count_18_io_out ? io_r_38_b : _GEN_7417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7419 = 9'h27 == r_count_18_io_out ? io_r_39_b : _GEN_7418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7420 = 9'h28 == r_count_18_io_out ? io_r_40_b : _GEN_7419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7421 = 9'h29 == r_count_18_io_out ? io_r_41_b : _GEN_7420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7422 = 9'h2a == r_count_18_io_out ? io_r_42_b : _GEN_7421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7423 = 9'h2b == r_count_18_io_out ? io_r_43_b : _GEN_7422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7424 = 9'h2c == r_count_18_io_out ? io_r_44_b : _GEN_7423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7425 = 9'h2d == r_count_18_io_out ? io_r_45_b : _GEN_7424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7426 = 9'h2e == r_count_18_io_out ? io_r_46_b : _GEN_7425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7427 = 9'h2f == r_count_18_io_out ? io_r_47_b : _GEN_7426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7428 = 9'h30 == r_count_18_io_out ? io_r_48_b : _GEN_7427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7429 = 9'h31 == r_count_18_io_out ? io_r_49_b : _GEN_7428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7430 = 9'h32 == r_count_18_io_out ? io_r_50_b : _GEN_7429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7431 = 9'h33 == r_count_18_io_out ? io_r_51_b : _GEN_7430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7432 = 9'h34 == r_count_18_io_out ? io_r_52_b : _GEN_7431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7433 = 9'h35 == r_count_18_io_out ? io_r_53_b : _GEN_7432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7434 = 9'h36 == r_count_18_io_out ? io_r_54_b : _GEN_7433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7435 = 9'h37 == r_count_18_io_out ? io_r_55_b : _GEN_7434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7436 = 9'h38 == r_count_18_io_out ? io_r_56_b : _GEN_7435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7437 = 9'h39 == r_count_18_io_out ? io_r_57_b : _GEN_7436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7438 = 9'h3a == r_count_18_io_out ? io_r_58_b : _GEN_7437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7439 = 9'h3b == r_count_18_io_out ? io_r_59_b : _GEN_7438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7440 = 9'h3c == r_count_18_io_out ? io_r_60_b : _GEN_7439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7441 = 9'h3d == r_count_18_io_out ? io_r_61_b : _GEN_7440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7442 = 9'h3e == r_count_18_io_out ? io_r_62_b : _GEN_7441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7443 = 9'h3f == r_count_18_io_out ? io_r_63_b : _GEN_7442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7444 = 9'h40 == r_count_18_io_out ? io_r_64_b : _GEN_7443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7445 = 9'h41 == r_count_18_io_out ? io_r_65_b : _GEN_7444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7446 = 9'h42 == r_count_18_io_out ? io_r_66_b : _GEN_7445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7447 = 9'h43 == r_count_18_io_out ? io_r_67_b : _GEN_7446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7448 = 9'h44 == r_count_18_io_out ? io_r_68_b : _GEN_7447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7449 = 9'h45 == r_count_18_io_out ? io_r_69_b : _GEN_7448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7450 = 9'h46 == r_count_18_io_out ? io_r_70_b : _GEN_7449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7451 = 9'h47 == r_count_18_io_out ? io_r_71_b : _GEN_7450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7452 = 9'h48 == r_count_18_io_out ? io_r_72_b : _GEN_7451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7453 = 9'h49 == r_count_18_io_out ? io_r_73_b : _GEN_7452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7454 = 9'h4a == r_count_18_io_out ? io_r_74_b : _GEN_7453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7455 = 9'h4b == r_count_18_io_out ? io_r_75_b : _GEN_7454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7456 = 9'h4c == r_count_18_io_out ? io_r_76_b : _GEN_7455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7457 = 9'h4d == r_count_18_io_out ? io_r_77_b : _GEN_7456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7458 = 9'h4e == r_count_18_io_out ? io_r_78_b : _GEN_7457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7459 = 9'h4f == r_count_18_io_out ? io_r_79_b : _GEN_7458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7460 = 9'h50 == r_count_18_io_out ? io_r_80_b : _GEN_7459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7461 = 9'h51 == r_count_18_io_out ? io_r_81_b : _GEN_7460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7462 = 9'h52 == r_count_18_io_out ? io_r_82_b : _GEN_7461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7463 = 9'h53 == r_count_18_io_out ? io_r_83_b : _GEN_7462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7464 = 9'h54 == r_count_18_io_out ? io_r_84_b : _GEN_7463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7465 = 9'h55 == r_count_18_io_out ? io_r_85_b : _GEN_7464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7466 = 9'h56 == r_count_18_io_out ? io_r_86_b : _GEN_7465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7467 = 9'h57 == r_count_18_io_out ? io_r_87_b : _GEN_7466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7468 = 9'h58 == r_count_18_io_out ? io_r_88_b : _GEN_7467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7469 = 9'h59 == r_count_18_io_out ? io_r_89_b : _GEN_7468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7470 = 9'h5a == r_count_18_io_out ? io_r_90_b : _GEN_7469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7471 = 9'h5b == r_count_18_io_out ? io_r_91_b : _GEN_7470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7472 = 9'h5c == r_count_18_io_out ? io_r_92_b : _GEN_7471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7473 = 9'h5d == r_count_18_io_out ? io_r_93_b : _GEN_7472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7474 = 9'h5e == r_count_18_io_out ? io_r_94_b : _GEN_7473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7475 = 9'h5f == r_count_18_io_out ? io_r_95_b : _GEN_7474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7476 = 9'h60 == r_count_18_io_out ? io_r_96_b : _GEN_7475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7477 = 9'h61 == r_count_18_io_out ? io_r_97_b : _GEN_7476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7478 = 9'h62 == r_count_18_io_out ? io_r_98_b : _GEN_7477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7479 = 9'h63 == r_count_18_io_out ? io_r_99_b : _GEN_7478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7480 = 9'h64 == r_count_18_io_out ? io_r_100_b : _GEN_7479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7481 = 9'h65 == r_count_18_io_out ? io_r_101_b : _GEN_7480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7482 = 9'h66 == r_count_18_io_out ? io_r_102_b : _GEN_7481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7483 = 9'h67 == r_count_18_io_out ? io_r_103_b : _GEN_7482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7484 = 9'h68 == r_count_18_io_out ? io_r_104_b : _GEN_7483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7485 = 9'h69 == r_count_18_io_out ? io_r_105_b : _GEN_7484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7486 = 9'h6a == r_count_18_io_out ? io_r_106_b : _GEN_7485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7487 = 9'h6b == r_count_18_io_out ? io_r_107_b : _GEN_7486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7488 = 9'h6c == r_count_18_io_out ? io_r_108_b : _GEN_7487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7489 = 9'h6d == r_count_18_io_out ? io_r_109_b : _GEN_7488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7490 = 9'h6e == r_count_18_io_out ? io_r_110_b : _GEN_7489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7491 = 9'h6f == r_count_18_io_out ? io_r_111_b : _GEN_7490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7492 = 9'h70 == r_count_18_io_out ? io_r_112_b : _GEN_7491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7493 = 9'h71 == r_count_18_io_out ? io_r_113_b : _GEN_7492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7494 = 9'h72 == r_count_18_io_out ? io_r_114_b : _GEN_7493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7495 = 9'h73 == r_count_18_io_out ? io_r_115_b : _GEN_7494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7496 = 9'h74 == r_count_18_io_out ? io_r_116_b : _GEN_7495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7497 = 9'h75 == r_count_18_io_out ? io_r_117_b : _GEN_7496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7498 = 9'h76 == r_count_18_io_out ? io_r_118_b : _GEN_7497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7499 = 9'h77 == r_count_18_io_out ? io_r_119_b : _GEN_7498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7500 = 9'h78 == r_count_18_io_out ? io_r_120_b : _GEN_7499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7501 = 9'h79 == r_count_18_io_out ? io_r_121_b : _GEN_7500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7502 = 9'h7a == r_count_18_io_out ? io_r_122_b : _GEN_7501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7503 = 9'h7b == r_count_18_io_out ? io_r_123_b : _GEN_7502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7504 = 9'h7c == r_count_18_io_out ? io_r_124_b : _GEN_7503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7505 = 9'h7d == r_count_18_io_out ? io_r_125_b : _GEN_7504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7506 = 9'h7e == r_count_18_io_out ? io_r_126_b : _GEN_7505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7507 = 9'h7f == r_count_18_io_out ? io_r_127_b : _GEN_7506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7508 = 9'h80 == r_count_18_io_out ? io_r_128_b : _GEN_7507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7509 = 9'h81 == r_count_18_io_out ? io_r_129_b : _GEN_7508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7510 = 9'h82 == r_count_18_io_out ? io_r_130_b : _GEN_7509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7511 = 9'h83 == r_count_18_io_out ? io_r_131_b : _GEN_7510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7512 = 9'h84 == r_count_18_io_out ? io_r_132_b : _GEN_7511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7513 = 9'h85 == r_count_18_io_out ? io_r_133_b : _GEN_7512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7514 = 9'h86 == r_count_18_io_out ? io_r_134_b : _GEN_7513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7515 = 9'h87 == r_count_18_io_out ? io_r_135_b : _GEN_7514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7516 = 9'h88 == r_count_18_io_out ? io_r_136_b : _GEN_7515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7517 = 9'h89 == r_count_18_io_out ? io_r_137_b : _GEN_7516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7518 = 9'h8a == r_count_18_io_out ? io_r_138_b : _GEN_7517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7519 = 9'h8b == r_count_18_io_out ? io_r_139_b : _GEN_7518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7520 = 9'h8c == r_count_18_io_out ? io_r_140_b : _GEN_7519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7521 = 9'h8d == r_count_18_io_out ? io_r_141_b : _GEN_7520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7522 = 9'h8e == r_count_18_io_out ? io_r_142_b : _GEN_7521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7523 = 9'h8f == r_count_18_io_out ? io_r_143_b : _GEN_7522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7524 = 9'h90 == r_count_18_io_out ? io_r_144_b : _GEN_7523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7525 = 9'h91 == r_count_18_io_out ? io_r_145_b : _GEN_7524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7526 = 9'h92 == r_count_18_io_out ? io_r_146_b : _GEN_7525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7527 = 9'h93 == r_count_18_io_out ? io_r_147_b : _GEN_7526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7528 = 9'h94 == r_count_18_io_out ? io_r_148_b : _GEN_7527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7529 = 9'h95 == r_count_18_io_out ? io_r_149_b : _GEN_7528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7530 = 9'h96 == r_count_18_io_out ? io_r_150_b : _GEN_7529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7531 = 9'h97 == r_count_18_io_out ? io_r_151_b : _GEN_7530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7532 = 9'h98 == r_count_18_io_out ? io_r_152_b : _GEN_7531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7533 = 9'h99 == r_count_18_io_out ? io_r_153_b : _GEN_7532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7534 = 9'h9a == r_count_18_io_out ? io_r_154_b : _GEN_7533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7535 = 9'h9b == r_count_18_io_out ? io_r_155_b : _GEN_7534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7536 = 9'h9c == r_count_18_io_out ? io_r_156_b : _GEN_7535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7537 = 9'h9d == r_count_18_io_out ? io_r_157_b : _GEN_7536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7538 = 9'h9e == r_count_18_io_out ? io_r_158_b : _GEN_7537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7539 = 9'h9f == r_count_18_io_out ? io_r_159_b : _GEN_7538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7540 = 9'ha0 == r_count_18_io_out ? io_r_160_b : _GEN_7539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7541 = 9'ha1 == r_count_18_io_out ? io_r_161_b : _GEN_7540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7542 = 9'ha2 == r_count_18_io_out ? io_r_162_b : _GEN_7541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7543 = 9'ha3 == r_count_18_io_out ? io_r_163_b : _GEN_7542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7544 = 9'ha4 == r_count_18_io_out ? io_r_164_b : _GEN_7543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7545 = 9'ha5 == r_count_18_io_out ? io_r_165_b : _GEN_7544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7546 = 9'ha6 == r_count_18_io_out ? io_r_166_b : _GEN_7545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7547 = 9'ha7 == r_count_18_io_out ? io_r_167_b : _GEN_7546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7548 = 9'ha8 == r_count_18_io_out ? io_r_168_b : _GEN_7547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7549 = 9'ha9 == r_count_18_io_out ? io_r_169_b : _GEN_7548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7550 = 9'haa == r_count_18_io_out ? io_r_170_b : _GEN_7549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7551 = 9'hab == r_count_18_io_out ? io_r_171_b : _GEN_7550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7552 = 9'hac == r_count_18_io_out ? io_r_172_b : _GEN_7551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7553 = 9'had == r_count_18_io_out ? io_r_173_b : _GEN_7552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7554 = 9'hae == r_count_18_io_out ? io_r_174_b : _GEN_7553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7555 = 9'haf == r_count_18_io_out ? io_r_175_b : _GEN_7554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7556 = 9'hb0 == r_count_18_io_out ? io_r_176_b : _GEN_7555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7557 = 9'hb1 == r_count_18_io_out ? io_r_177_b : _GEN_7556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7558 = 9'hb2 == r_count_18_io_out ? io_r_178_b : _GEN_7557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7559 = 9'hb3 == r_count_18_io_out ? io_r_179_b : _GEN_7558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7560 = 9'hb4 == r_count_18_io_out ? io_r_180_b : _GEN_7559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7561 = 9'hb5 == r_count_18_io_out ? io_r_181_b : _GEN_7560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7562 = 9'hb6 == r_count_18_io_out ? io_r_182_b : _GEN_7561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7563 = 9'hb7 == r_count_18_io_out ? io_r_183_b : _GEN_7562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7564 = 9'hb8 == r_count_18_io_out ? io_r_184_b : _GEN_7563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7565 = 9'hb9 == r_count_18_io_out ? io_r_185_b : _GEN_7564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7566 = 9'hba == r_count_18_io_out ? io_r_186_b : _GEN_7565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7567 = 9'hbb == r_count_18_io_out ? io_r_187_b : _GEN_7566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7568 = 9'hbc == r_count_18_io_out ? io_r_188_b : _GEN_7567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7569 = 9'hbd == r_count_18_io_out ? io_r_189_b : _GEN_7568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7570 = 9'hbe == r_count_18_io_out ? io_r_190_b : _GEN_7569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7571 = 9'hbf == r_count_18_io_out ? io_r_191_b : _GEN_7570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7572 = 9'hc0 == r_count_18_io_out ? io_r_192_b : _GEN_7571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7573 = 9'hc1 == r_count_18_io_out ? io_r_193_b : _GEN_7572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7574 = 9'hc2 == r_count_18_io_out ? io_r_194_b : _GEN_7573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7575 = 9'hc3 == r_count_18_io_out ? io_r_195_b : _GEN_7574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7576 = 9'hc4 == r_count_18_io_out ? io_r_196_b : _GEN_7575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7577 = 9'hc5 == r_count_18_io_out ? io_r_197_b : _GEN_7576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7578 = 9'hc6 == r_count_18_io_out ? io_r_198_b : _GEN_7577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7579 = 9'hc7 == r_count_18_io_out ? io_r_199_b : _GEN_7578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7580 = 9'hc8 == r_count_18_io_out ? io_r_200_b : _GEN_7579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7581 = 9'hc9 == r_count_18_io_out ? io_r_201_b : _GEN_7580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7582 = 9'hca == r_count_18_io_out ? io_r_202_b : _GEN_7581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7583 = 9'hcb == r_count_18_io_out ? io_r_203_b : _GEN_7582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7584 = 9'hcc == r_count_18_io_out ? io_r_204_b : _GEN_7583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7585 = 9'hcd == r_count_18_io_out ? io_r_205_b : _GEN_7584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7586 = 9'hce == r_count_18_io_out ? io_r_206_b : _GEN_7585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7587 = 9'hcf == r_count_18_io_out ? io_r_207_b : _GEN_7586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7588 = 9'hd0 == r_count_18_io_out ? io_r_208_b : _GEN_7587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7589 = 9'hd1 == r_count_18_io_out ? io_r_209_b : _GEN_7588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7590 = 9'hd2 == r_count_18_io_out ? io_r_210_b : _GEN_7589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7591 = 9'hd3 == r_count_18_io_out ? io_r_211_b : _GEN_7590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7592 = 9'hd4 == r_count_18_io_out ? io_r_212_b : _GEN_7591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7593 = 9'hd5 == r_count_18_io_out ? io_r_213_b : _GEN_7592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7594 = 9'hd6 == r_count_18_io_out ? io_r_214_b : _GEN_7593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7595 = 9'hd7 == r_count_18_io_out ? io_r_215_b : _GEN_7594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7596 = 9'hd8 == r_count_18_io_out ? io_r_216_b : _GEN_7595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7597 = 9'hd9 == r_count_18_io_out ? io_r_217_b : _GEN_7596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7598 = 9'hda == r_count_18_io_out ? io_r_218_b : _GEN_7597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7599 = 9'hdb == r_count_18_io_out ? io_r_219_b : _GEN_7598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7600 = 9'hdc == r_count_18_io_out ? io_r_220_b : _GEN_7599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7601 = 9'hdd == r_count_18_io_out ? io_r_221_b : _GEN_7600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7602 = 9'hde == r_count_18_io_out ? io_r_222_b : _GEN_7601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7603 = 9'hdf == r_count_18_io_out ? io_r_223_b : _GEN_7602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7604 = 9'he0 == r_count_18_io_out ? io_r_224_b : _GEN_7603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7605 = 9'he1 == r_count_18_io_out ? io_r_225_b : _GEN_7604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7606 = 9'he2 == r_count_18_io_out ? io_r_226_b : _GEN_7605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7607 = 9'he3 == r_count_18_io_out ? io_r_227_b : _GEN_7606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7608 = 9'he4 == r_count_18_io_out ? io_r_228_b : _GEN_7607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7609 = 9'he5 == r_count_18_io_out ? io_r_229_b : _GEN_7608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7610 = 9'he6 == r_count_18_io_out ? io_r_230_b : _GEN_7609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7611 = 9'he7 == r_count_18_io_out ? io_r_231_b : _GEN_7610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7612 = 9'he8 == r_count_18_io_out ? io_r_232_b : _GEN_7611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7613 = 9'he9 == r_count_18_io_out ? io_r_233_b : _GEN_7612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7614 = 9'hea == r_count_18_io_out ? io_r_234_b : _GEN_7613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7615 = 9'heb == r_count_18_io_out ? io_r_235_b : _GEN_7614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7616 = 9'hec == r_count_18_io_out ? io_r_236_b : _GEN_7615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7617 = 9'hed == r_count_18_io_out ? io_r_237_b : _GEN_7616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7618 = 9'hee == r_count_18_io_out ? io_r_238_b : _GEN_7617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7619 = 9'hef == r_count_18_io_out ? io_r_239_b : _GEN_7618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7620 = 9'hf0 == r_count_18_io_out ? io_r_240_b : _GEN_7619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7621 = 9'hf1 == r_count_18_io_out ? io_r_241_b : _GEN_7620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7622 = 9'hf2 == r_count_18_io_out ? io_r_242_b : _GEN_7621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7623 = 9'hf3 == r_count_18_io_out ? io_r_243_b : _GEN_7622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7624 = 9'hf4 == r_count_18_io_out ? io_r_244_b : _GEN_7623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7625 = 9'hf5 == r_count_18_io_out ? io_r_245_b : _GEN_7624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7626 = 9'hf6 == r_count_18_io_out ? io_r_246_b : _GEN_7625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7627 = 9'hf7 == r_count_18_io_out ? io_r_247_b : _GEN_7626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7628 = 9'hf8 == r_count_18_io_out ? io_r_248_b : _GEN_7627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7629 = 9'hf9 == r_count_18_io_out ? io_r_249_b : _GEN_7628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7630 = 9'hfa == r_count_18_io_out ? io_r_250_b : _GEN_7629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7631 = 9'hfb == r_count_18_io_out ? io_r_251_b : _GEN_7630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7632 = 9'hfc == r_count_18_io_out ? io_r_252_b : _GEN_7631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7633 = 9'hfd == r_count_18_io_out ? io_r_253_b : _GEN_7632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7634 = 9'hfe == r_count_18_io_out ? io_r_254_b : _GEN_7633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7635 = 9'hff == r_count_18_io_out ? io_r_255_b : _GEN_7634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7636 = 9'h100 == r_count_18_io_out ? io_r_256_b : _GEN_7635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7637 = 9'h101 == r_count_18_io_out ? io_r_257_b : _GEN_7636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7638 = 9'h102 == r_count_18_io_out ? io_r_258_b : _GEN_7637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7639 = 9'h103 == r_count_18_io_out ? io_r_259_b : _GEN_7638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7640 = 9'h104 == r_count_18_io_out ? io_r_260_b : _GEN_7639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7641 = 9'h105 == r_count_18_io_out ? io_r_261_b : _GEN_7640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7642 = 9'h106 == r_count_18_io_out ? io_r_262_b : _GEN_7641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7643 = 9'h107 == r_count_18_io_out ? io_r_263_b : _GEN_7642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7644 = 9'h108 == r_count_18_io_out ? io_r_264_b : _GEN_7643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7645 = 9'h109 == r_count_18_io_out ? io_r_265_b : _GEN_7644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7646 = 9'h10a == r_count_18_io_out ? io_r_266_b : _GEN_7645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7647 = 9'h10b == r_count_18_io_out ? io_r_267_b : _GEN_7646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7648 = 9'h10c == r_count_18_io_out ? io_r_268_b : _GEN_7647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7649 = 9'h10d == r_count_18_io_out ? io_r_269_b : _GEN_7648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7650 = 9'h10e == r_count_18_io_out ? io_r_270_b : _GEN_7649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7651 = 9'h10f == r_count_18_io_out ? io_r_271_b : _GEN_7650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7652 = 9'h110 == r_count_18_io_out ? io_r_272_b : _GEN_7651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7653 = 9'h111 == r_count_18_io_out ? io_r_273_b : _GEN_7652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7654 = 9'h112 == r_count_18_io_out ? io_r_274_b : _GEN_7653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7655 = 9'h113 == r_count_18_io_out ? io_r_275_b : _GEN_7654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7656 = 9'h114 == r_count_18_io_out ? io_r_276_b : _GEN_7655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7657 = 9'h115 == r_count_18_io_out ? io_r_277_b : _GEN_7656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7658 = 9'h116 == r_count_18_io_out ? io_r_278_b : _GEN_7657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7659 = 9'h117 == r_count_18_io_out ? io_r_279_b : _GEN_7658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7660 = 9'h118 == r_count_18_io_out ? io_r_280_b : _GEN_7659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7661 = 9'h119 == r_count_18_io_out ? io_r_281_b : _GEN_7660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7662 = 9'h11a == r_count_18_io_out ? io_r_282_b : _GEN_7661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7663 = 9'h11b == r_count_18_io_out ? io_r_283_b : _GEN_7662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7664 = 9'h11c == r_count_18_io_out ? io_r_284_b : _GEN_7663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7665 = 9'h11d == r_count_18_io_out ? io_r_285_b : _GEN_7664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7666 = 9'h11e == r_count_18_io_out ? io_r_286_b : _GEN_7665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7667 = 9'h11f == r_count_18_io_out ? io_r_287_b : _GEN_7666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7668 = 9'h120 == r_count_18_io_out ? io_r_288_b : _GEN_7667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7669 = 9'h121 == r_count_18_io_out ? io_r_289_b : _GEN_7668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7670 = 9'h122 == r_count_18_io_out ? io_r_290_b : _GEN_7669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7671 = 9'h123 == r_count_18_io_out ? io_r_291_b : _GEN_7670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7672 = 9'h124 == r_count_18_io_out ? io_r_292_b : _GEN_7671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7673 = 9'h125 == r_count_18_io_out ? io_r_293_b : _GEN_7672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7674 = 9'h126 == r_count_18_io_out ? io_r_294_b : _GEN_7673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7675 = 9'h127 == r_count_18_io_out ? io_r_295_b : _GEN_7674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7676 = 9'h128 == r_count_18_io_out ? io_r_296_b : _GEN_7675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7677 = 9'h129 == r_count_18_io_out ? io_r_297_b : _GEN_7676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7678 = 9'h12a == r_count_18_io_out ? io_r_298_b : _GEN_7677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7679 = 9'h12b == r_count_18_io_out ? io_r_299_b : _GEN_7678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7680 = 9'h12c == r_count_18_io_out ? io_r_300_b : _GEN_7679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7681 = 9'h12d == r_count_18_io_out ? io_r_301_b : _GEN_7680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7682 = 9'h12e == r_count_18_io_out ? io_r_302_b : _GEN_7681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7683 = 9'h12f == r_count_18_io_out ? io_r_303_b : _GEN_7682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7684 = 9'h130 == r_count_18_io_out ? io_r_304_b : _GEN_7683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7685 = 9'h131 == r_count_18_io_out ? io_r_305_b : _GEN_7684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7686 = 9'h132 == r_count_18_io_out ? io_r_306_b : _GEN_7685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7687 = 9'h133 == r_count_18_io_out ? io_r_307_b : _GEN_7686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7688 = 9'h134 == r_count_18_io_out ? io_r_308_b : _GEN_7687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7689 = 9'h135 == r_count_18_io_out ? io_r_309_b : _GEN_7688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7690 = 9'h136 == r_count_18_io_out ? io_r_310_b : _GEN_7689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7691 = 9'h137 == r_count_18_io_out ? io_r_311_b : _GEN_7690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7692 = 9'h138 == r_count_18_io_out ? io_r_312_b : _GEN_7691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7693 = 9'h139 == r_count_18_io_out ? io_r_313_b : _GEN_7692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7694 = 9'h13a == r_count_18_io_out ? io_r_314_b : _GEN_7693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7695 = 9'h13b == r_count_18_io_out ? io_r_315_b : _GEN_7694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7696 = 9'h13c == r_count_18_io_out ? io_r_316_b : _GEN_7695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7697 = 9'h13d == r_count_18_io_out ? io_r_317_b : _GEN_7696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7698 = 9'h13e == r_count_18_io_out ? io_r_318_b : _GEN_7697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7699 = 9'h13f == r_count_18_io_out ? io_r_319_b : _GEN_7698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7700 = 9'h140 == r_count_18_io_out ? io_r_320_b : _GEN_7699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7701 = 9'h141 == r_count_18_io_out ? io_r_321_b : _GEN_7700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7702 = 9'h142 == r_count_18_io_out ? io_r_322_b : _GEN_7701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7703 = 9'h143 == r_count_18_io_out ? io_r_323_b : _GEN_7702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7704 = 9'h144 == r_count_18_io_out ? io_r_324_b : _GEN_7703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7705 = 9'h145 == r_count_18_io_out ? io_r_325_b : _GEN_7704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7706 = 9'h146 == r_count_18_io_out ? io_r_326_b : _GEN_7705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7707 = 9'h147 == r_count_18_io_out ? io_r_327_b : _GEN_7706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7708 = 9'h148 == r_count_18_io_out ? io_r_328_b : _GEN_7707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7709 = 9'h149 == r_count_18_io_out ? io_r_329_b : _GEN_7708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7710 = 9'h14a == r_count_18_io_out ? io_r_330_b : _GEN_7709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7711 = 9'h14b == r_count_18_io_out ? io_r_331_b : _GEN_7710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7712 = 9'h14c == r_count_18_io_out ? io_r_332_b : _GEN_7711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7713 = 9'h14d == r_count_18_io_out ? io_r_333_b : _GEN_7712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7714 = 9'h14e == r_count_18_io_out ? io_r_334_b : _GEN_7713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7715 = 9'h14f == r_count_18_io_out ? io_r_335_b : _GEN_7714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7716 = 9'h150 == r_count_18_io_out ? io_r_336_b : _GEN_7715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7717 = 9'h151 == r_count_18_io_out ? io_r_337_b : _GEN_7716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7718 = 9'h152 == r_count_18_io_out ? io_r_338_b : _GEN_7717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7719 = 9'h153 == r_count_18_io_out ? io_r_339_b : _GEN_7718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7720 = 9'h154 == r_count_18_io_out ? io_r_340_b : _GEN_7719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7721 = 9'h155 == r_count_18_io_out ? io_r_341_b : _GEN_7720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7722 = 9'h156 == r_count_18_io_out ? io_r_342_b : _GEN_7721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7723 = 9'h157 == r_count_18_io_out ? io_r_343_b : _GEN_7722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7724 = 9'h158 == r_count_18_io_out ? io_r_344_b : _GEN_7723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7725 = 9'h159 == r_count_18_io_out ? io_r_345_b : _GEN_7724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7726 = 9'h15a == r_count_18_io_out ? io_r_346_b : _GEN_7725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7727 = 9'h15b == r_count_18_io_out ? io_r_347_b : _GEN_7726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7728 = 9'h15c == r_count_18_io_out ? io_r_348_b : _GEN_7727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7729 = 9'h15d == r_count_18_io_out ? io_r_349_b : _GEN_7728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7730 = 9'h15e == r_count_18_io_out ? io_r_350_b : _GEN_7729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7731 = 9'h15f == r_count_18_io_out ? io_r_351_b : _GEN_7730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7732 = 9'h160 == r_count_18_io_out ? io_r_352_b : _GEN_7731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7733 = 9'h161 == r_count_18_io_out ? io_r_353_b : _GEN_7732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7734 = 9'h162 == r_count_18_io_out ? io_r_354_b : _GEN_7733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7735 = 9'h163 == r_count_18_io_out ? io_r_355_b : _GEN_7734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7736 = 9'h164 == r_count_18_io_out ? io_r_356_b : _GEN_7735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7737 = 9'h165 == r_count_18_io_out ? io_r_357_b : _GEN_7736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7738 = 9'h166 == r_count_18_io_out ? io_r_358_b : _GEN_7737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7739 = 9'h167 == r_count_18_io_out ? io_r_359_b : _GEN_7738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7740 = 9'h168 == r_count_18_io_out ? io_r_360_b : _GEN_7739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7741 = 9'h169 == r_count_18_io_out ? io_r_361_b : _GEN_7740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7742 = 9'h16a == r_count_18_io_out ? io_r_362_b : _GEN_7741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7743 = 9'h16b == r_count_18_io_out ? io_r_363_b : _GEN_7742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7744 = 9'h16c == r_count_18_io_out ? io_r_364_b : _GEN_7743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7745 = 9'h16d == r_count_18_io_out ? io_r_365_b : _GEN_7744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7746 = 9'h16e == r_count_18_io_out ? io_r_366_b : _GEN_7745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7747 = 9'h16f == r_count_18_io_out ? io_r_367_b : _GEN_7746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7748 = 9'h170 == r_count_18_io_out ? io_r_368_b : _GEN_7747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7749 = 9'h171 == r_count_18_io_out ? io_r_369_b : _GEN_7748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7750 = 9'h172 == r_count_18_io_out ? io_r_370_b : _GEN_7749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7751 = 9'h173 == r_count_18_io_out ? io_r_371_b : _GEN_7750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7752 = 9'h174 == r_count_18_io_out ? io_r_372_b : _GEN_7751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7753 = 9'h175 == r_count_18_io_out ? io_r_373_b : _GEN_7752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7754 = 9'h176 == r_count_18_io_out ? io_r_374_b : _GEN_7753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7755 = 9'h177 == r_count_18_io_out ? io_r_375_b : _GEN_7754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7756 = 9'h178 == r_count_18_io_out ? io_r_376_b : _GEN_7755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7757 = 9'h179 == r_count_18_io_out ? io_r_377_b : _GEN_7756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7758 = 9'h17a == r_count_18_io_out ? io_r_378_b : _GEN_7757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7759 = 9'h17b == r_count_18_io_out ? io_r_379_b : _GEN_7758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7760 = 9'h17c == r_count_18_io_out ? io_r_380_b : _GEN_7759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7761 = 9'h17d == r_count_18_io_out ? io_r_381_b : _GEN_7760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7762 = 9'h17e == r_count_18_io_out ? io_r_382_b : _GEN_7761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7763 = 9'h17f == r_count_18_io_out ? io_r_383_b : _GEN_7762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7764 = 9'h180 == r_count_18_io_out ? io_r_384_b : _GEN_7763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7765 = 9'h181 == r_count_18_io_out ? io_r_385_b : _GEN_7764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7766 = 9'h182 == r_count_18_io_out ? io_r_386_b : _GEN_7765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7767 = 9'h183 == r_count_18_io_out ? io_r_387_b : _GEN_7766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7768 = 9'h184 == r_count_18_io_out ? io_r_388_b : _GEN_7767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7769 = 9'h185 == r_count_18_io_out ? io_r_389_b : _GEN_7768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7770 = 9'h186 == r_count_18_io_out ? io_r_390_b : _GEN_7769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7771 = 9'h187 == r_count_18_io_out ? io_r_391_b : _GEN_7770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7772 = 9'h188 == r_count_18_io_out ? io_r_392_b : _GEN_7771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7773 = 9'h189 == r_count_18_io_out ? io_r_393_b : _GEN_7772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7774 = 9'h18a == r_count_18_io_out ? io_r_394_b : _GEN_7773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7775 = 9'h18b == r_count_18_io_out ? io_r_395_b : _GEN_7774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7776 = 9'h18c == r_count_18_io_out ? io_r_396_b : _GEN_7775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7777 = 9'h18d == r_count_18_io_out ? io_r_397_b : _GEN_7776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7778 = 9'h18e == r_count_18_io_out ? io_r_398_b : _GEN_7777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7781 = 9'h1 == r_count_19_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7782 = 9'h2 == r_count_19_io_out ? io_r_2_b : _GEN_7781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7783 = 9'h3 == r_count_19_io_out ? io_r_3_b : _GEN_7782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7784 = 9'h4 == r_count_19_io_out ? io_r_4_b : _GEN_7783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7785 = 9'h5 == r_count_19_io_out ? io_r_5_b : _GEN_7784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7786 = 9'h6 == r_count_19_io_out ? io_r_6_b : _GEN_7785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7787 = 9'h7 == r_count_19_io_out ? io_r_7_b : _GEN_7786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7788 = 9'h8 == r_count_19_io_out ? io_r_8_b : _GEN_7787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7789 = 9'h9 == r_count_19_io_out ? io_r_9_b : _GEN_7788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7790 = 9'ha == r_count_19_io_out ? io_r_10_b : _GEN_7789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7791 = 9'hb == r_count_19_io_out ? io_r_11_b : _GEN_7790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7792 = 9'hc == r_count_19_io_out ? io_r_12_b : _GEN_7791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7793 = 9'hd == r_count_19_io_out ? io_r_13_b : _GEN_7792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7794 = 9'he == r_count_19_io_out ? io_r_14_b : _GEN_7793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7795 = 9'hf == r_count_19_io_out ? io_r_15_b : _GEN_7794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7796 = 9'h10 == r_count_19_io_out ? io_r_16_b : _GEN_7795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7797 = 9'h11 == r_count_19_io_out ? io_r_17_b : _GEN_7796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7798 = 9'h12 == r_count_19_io_out ? io_r_18_b : _GEN_7797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7799 = 9'h13 == r_count_19_io_out ? io_r_19_b : _GEN_7798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7800 = 9'h14 == r_count_19_io_out ? io_r_20_b : _GEN_7799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7801 = 9'h15 == r_count_19_io_out ? io_r_21_b : _GEN_7800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7802 = 9'h16 == r_count_19_io_out ? io_r_22_b : _GEN_7801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7803 = 9'h17 == r_count_19_io_out ? io_r_23_b : _GEN_7802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7804 = 9'h18 == r_count_19_io_out ? io_r_24_b : _GEN_7803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7805 = 9'h19 == r_count_19_io_out ? io_r_25_b : _GEN_7804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7806 = 9'h1a == r_count_19_io_out ? io_r_26_b : _GEN_7805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7807 = 9'h1b == r_count_19_io_out ? io_r_27_b : _GEN_7806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7808 = 9'h1c == r_count_19_io_out ? io_r_28_b : _GEN_7807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7809 = 9'h1d == r_count_19_io_out ? io_r_29_b : _GEN_7808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7810 = 9'h1e == r_count_19_io_out ? io_r_30_b : _GEN_7809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7811 = 9'h1f == r_count_19_io_out ? io_r_31_b : _GEN_7810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7812 = 9'h20 == r_count_19_io_out ? io_r_32_b : _GEN_7811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7813 = 9'h21 == r_count_19_io_out ? io_r_33_b : _GEN_7812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7814 = 9'h22 == r_count_19_io_out ? io_r_34_b : _GEN_7813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7815 = 9'h23 == r_count_19_io_out ? io_r_35_b : _GEN_7814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7816 = 9'h24 == r_count_19_io_out ? io_r_36_b : _GEN_7815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7817 = 9'h25 == r_count_19_io_out ? io_r_37_b : _GEN_7816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7818 = 9'h26 == r_count_19_io_out ? io_r_38_b : _GEN_7817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7819 = 9'h27 == r_count_19_io_out ? io_r_39_b : _GEN_7818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7820 = 9'h28 == r_count_19_io_out ? io_r_40_b : _GEN_7819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7821 = 9'h29 == r_count_19_io_out ? io_r_41_b : _GEN_7820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7822 = 9'h2a == r_count_19_io_out ? io_r_42_b : _GEN_7821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7823 = 9'h2b == r_count_19_io_out ? io_r_43_b : _GEN_7822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7824 = 9'h2c == r_count_19_io_out ? io_r_44_b : _GEN_7823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7825 = 9'h2d == r_count_19_io_out ? io_r_45_b : _GEN_7824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7826 = 9'h2e == r_count_19_io_out ? io_r_46_b : _GEN_7825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7827 = 9'h2f == r_count_19_io_out ? io_r_47_b : _GEN_7826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7828 = 9'h30 == r_count_19_io_out ? io_r_48_b : _GEN_7827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7829 = 9'h31 == r_count_19_io_out ? io_r_49_b : _GEN_7828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7830 = 9'h32 == r_count_19_io_out ? io_r_50_b : _GEN_7829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7831 = 9'h33 == r_count_19_io_out ? io_r_51_b : _GEN_7830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7832 = 9'h34 == r_count_19_io_out ? io_r_52_b : _GEN_7831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7833 = 9'h35 == r_count_19_io_out ? io_r_53_b : _GEN_7832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7834 = 9'h36 == r_count_19_io_out ? io_r_54_b : _GEN_7833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7835 = 9'h37 == r_count_19_io_out ? io_r_55_b : _GEN_7834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7836 = 9'h38 == r_count_19_io_out ? io_r_56_b : _GEN_7835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7837 = 9'h39 == r_count_19_io_out ? io_r_57_b : _GEN_7836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7838 = 9'h3a == r_count_19_io_out ? io_r_58_b : _GEN_7837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7839 = 9'h3b == r_count_19_io_out ? io_r_59_b : _GEN_7838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7840 = 9'h3c == r_count_19_io_out ? io_r_60_b : _GEN_7839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7841 = 9'h3d == r_count_19_io_out ? io_r_61_b : _GEN_7840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7842 = 9'h3e == r_count_19_io_out ? io_r_62_b : _GEN_7841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7843 = 9'h3f == r_count_19_io_out ? io_r_63_b : _GEN_7842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7844 = 9'h40 == r_count_19_io_out ? io_r_64_b : _GEN_7843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7845 = 9'h41 == r_count_19_io_out ? io_r_65_b : _GEN_7844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7846 = 9'h42 == r_count_19_io_out ? io_r_66_b : _GEN_7845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7847 = 9'h43 == r_count_19_io_out ? io_r_67_b : _GEN_7846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7848 = 9'h44 == r_count_19_io_out ? io_r_68_b : _GEN_7847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7849 = 9'h45 == r_count_19_io_out ? io_r_69_b : _GEN_7848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7850 = 9'h46 == r_count_19_io_out ? io_r_70_b : _GEN_7849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7851 = 9'h47 == r_count_19_io_out ? io_r_71_b : _GEN_7850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7852 = 9'h48 == r_count_19_io_out ? io_r_72_b : _GEN_7851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7853 = 9'h49 == r_count_19_io_out ? io_r_73_b : _GEN_7852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7854 = 9'h4a == r_count_19_io_out ? io_r_74_b : _GEN_7853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7855 = 9'h4b == r_count_19_io_out ? io_r_75_b : _GEN_7854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7856 = 9'h4c == r_count_19_io_out ? io_r_76_b : _GEN_7855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7857 = 9'h4d == r_count_19_io_out ? io_r_77_b : _GEN_7856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7858 = 9'h4e == r_count_19_io_out ? io_r_78_b : _GEN_7857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7859 = 9'h4f == r_count_19_io_out ? io_r_79_b : _GEN_7858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7860 = 9'h50 == r_count_19_io_out ? io_r_80_b : _GEN_7859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7861 = 9'h51 == r_count_19_io_out ? io_r_81_b : _GEN_7860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7862 = 9'h52 == r_count_19_io_out ? io_r_82_b : _GEN_7861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7863 = 9'h53 == r_count_19_io_out ? io_r_83_b : _GEN_7862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7864 = 9'h54 == r_count_19_io_out ? io_r_84_b : _GEN_7863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7865 = 9'h55 == r_count_19_io_out ? io_r_85_b : _GEN_7864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7866 = 9'h56 == r_count_19_io_out ? io_r_86_b : _GEN_7865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7867 = 9'h57 == r_count_19_io_out ? io_r_87_b : _GEN_7866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7868 = 9'h58 == r_count_19_io_out ? io_r_88_b : _GEN_7867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7869 = 9'h59 == r_count_19_io_out ? io_r_89_b : _GEN_7868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7870 = 9'h5a == r_count_19_io_out ? io_r_90_b : _GEN_7869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7871 = 9'h5b == r_count_19_io_out ? io_r_91_b : _GEN_7870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7872 = 9'h5c == r_count_19_io_out ? io_r_92_b : _GEN_7871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7873 = 9'h5d == r_count_19_io_out ? io_r_93_b : _GEN_7872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7874 = 9'h5e == r_count_19_io_out ? io_r_94_b : _GEN_7873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7875 = 9'h5f == r_count_19_io_out ? io_r_95_b : _GEN_7874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7876 = 9'h60 == r_count_19_io_out ? io_r_96_b : _GEN_7875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7877 = 9'h61 == r_count_19_io_out ? io_r_97_b : _GEN_7876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7878 = 9'h62 == r_count_19_io_out ? io_r_98_b : _GEN_7877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7879 = 9'h63 == r_count_19_io_out ? io_r_99_b : _GEN_7878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7880 = 9'h64 == r_count_19_io_out ? io_r_100_b : _GEN_7879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7881 = 9'h65 == r_count_19_io_out ? io_r_101_b : _GEN_7880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7882 = 9'h66 == r_count_19_io_out ? io_r_102_b : _GEN_7881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7883 = 9'h67 == r_count_19_io_out ? io_r_103_b : _GEN_7882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7884 = 9'h68 == r_count_19_io_out ? io_r_104_b : _GEN_7883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7885 = 9'h69 == r_count_19_io_out ? io_r_105_b : _GEN_7884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7886 = 9'h6a == r_count_19_io_out ? io_r_106_b : _GEN_7885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7887 = 9'h6b == r_count_19_io_out ? io_r_107_b : _GEN_7886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7888 = 9'h6c == r_count_19_io_out ? io_r_108_b : _GEN_7887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7889 = 9'h6d == r_count_19_io_out ? io_r_109_b : _GEN_7888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7890 = 9'h6e == r_count_19_io_out ? io_r_110_b : _GEN_7889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7891 = 9'h6f == r_count_19_io_out ? io_r_111_b : _GEN_7890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7892 = 9'h70 == r_count_19_io_out ? io_r_112_b : _GEN_7891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7893 = 9'h71 == r_count_19_io_out ? io_r_113_b : _GEN_7892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7894 = 9'h72 == r_count_19_io_out ? io_r_114_b : _GEN_7893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7895 = 9'h73 == r_count_19_io_out ? io_r_115_b : _GEN_7894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7896 = 9'h74 == r_count_19_io_out ? io_r_116_b : _GEN_7895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7897 = 9'h75 == r_count_19_io_out ? io_r_117_b : _GEN_7896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7898 = 9'h76 == r_count_19_io_out ? io_r_118_b : _GEN_7897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7899 = 9'h77 == r_count_19_io_out ? io_r_119_b : _GEN_7898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7900 = 9'h78 == r_count_19_io_out ? io_r_120_b : _GEN_7899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7901 = 9'h79 == r_count_19_io_out ? io_r_121_b : _GEN_7900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7902 = 9'h7a == r_count_19_io_out ? io_r_122_b : _GEN_7901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7903 = 9'h7b == r_count_19_io_out ? io_r_123_b : _GEN_7902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7904 = 9'h7c == r_count_19_io_out ? io_r_124_b : _GEN_7903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7905 = 9'h7d == r_count_19_io_out ? io_r_125_b : _GEN_7904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7906 = 9'h7e == r_count_19_io_out ? io_r_126_b : _GEN_7905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7907 = 9'h7f == r_count_19_io_out ? io_r_127_b : _GEN_7906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7908 = 9'h80 == r_count_19_io_out ? io_r_128_b : _GEN_7907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7909 = 9'h81 == r_count_19_io_out ? io_r_129_b : _GEN_7908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7910 = 9'h82 == r_count_19_io_out ? io_r_130_b : _GEN_7909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7911 = 9'h83 == r_count_19_io_out ? io_r_131_b : _GEN_7910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7912 = 9'h84 == r_count_19_io_out ? io_r_132_b : _GEN_7911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7913 = 9'h85 == r_count_19_io_out ? io_r_133_b : _GEN_7912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7914 = 9'h86 == r_count_19_io_out ? io_r_134_b : _GEN_7913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7915 = 9'h87 == r_count_19_io_out ? io_r_135_b : _GEN_7914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7916 = 9'h88 == r_count_19_io_out ? io_r_136_b : _GEN_7915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7917 = 9'h89 == r_count_19_io_out ? io_r_137_b : _GEN_7916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7918 = 9'h8a == r_count_19_io_out ? io_r_138_b : _GEN_7917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7919 = 9'h8b == r_count_19_io_out ? io_r_139_b : _GEN_7918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7920 = 9'h8c == r_count_19_io_out ? io_r_140_b : _GEN_7919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7921 = 9'h8d == r_count_19_io_out ? io_r_141_b : _GEN_7920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7922 = 9'h8e == r_count_19_io_out ? io_r_142_b : _GEN_7921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7923 = 9'h8f == r_count_19_io_out ? io_r_143_b : _GEN_7922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7924 = 9'h90 == r_count_19_io_out ? io_r_144_b : _GEN_7923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7925 = 9'h91 == r_count_19_io_out ? io_r_145_b : _GEN_7924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7926 = 9'h92 == r_count_19_io_out ? io_r_146_b : _GEN_7925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7927 = 9'h93 == r_count_19_io_out ? io_r_147_b : _GEN_7926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7928 = 9'h94 == r_count_19_io_out ? io_r_148_b : _GEN_7927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7929 = 9'h95 == r_count_19_io_out ? io_r_149_b : _GEN_7928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7930 = 9'h96 == r_count_19_io_out ? io_r_150_b : _GEN_7929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7931 = 9'h97 == r_count_19_io_out ? io_r_151_b : _GEN_7930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7932 = 9'h98 == r_count_19_io_out ? io_r_152_b : _GEN_7931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7933 = 9'h99 == r_count_19_io_out ? io_r_153_b : _GEN_7932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7934 = 9'h9a == r_count_19_io_out ? io_r_154_b : _GEN_7933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7935 = 9'h9b == r_count_19_io_out ? io_r_155_b : _GEN_7934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7936 = 9'h9c == r_count_19_io_out ? io_r_156_b : _GEN_7935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7937 = 9'h9d == r_count_19_io_out ? io_r_157_b : _GEN_7936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7938 = 9'h9e == r_count_19_io_out ? io_r_158_b : _GEN_7937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7939 = 9'h9f == r_count_19_io_out ? io_r_159_b : _GEN_7938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7940 = 9'ha0 == r_count_19_io_out ? io_r_160_b : _GEN_7939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7941 = 9'ha1 == r_count_19_io_out ? io_r_161_b : _GEN_7940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7942 = 9'ha2 == r_count_19_io_out ? io_r_162_b : _GEN_7941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7943 = 9'ha3 == r_count_19_io_out ? io_r_163_b : _GEN_7942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7944 = 9'ha4 == r_count_19_io_out ? io_r_164_b : _GEN_7943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7945 = 9'ha5 == r_count_19_io_out ? io_r_165_b : _GEN_7944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7946 = 9'ha6 == r_count_19_io_out ? io_r_166_b : _GEN_7945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7947 = 9'ha7 == r_count_19_io_out ? io_r_167_b : _GEN_7946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7948 = 9'ha8 == r_count_19_io_out ? io_r_168_b : _GEN_7947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7949 = 9'ha9 == r_count_19_io_out ? io_r_169_b : _GEN_7948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7950 = 9'haa == r_count_19_io_out ? io_r_170_b : _GEN_7949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7951 = 9'hab == r_count_19_io_out ? io_r_171_b : _GEN_7950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7952 = 9'hac == r_count_19_io_out ? io_r_172_b : _GEN_7951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7953 = 9'had == r_count_19_io_out ? io_r_173_b : _GEN_7952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7954 = 9'hae == r_count_19_io_out ? io_r_174_b : _GEN_7953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7955 = 9'haf == r_count_19_io_out ? io_r_175_b : _GEN_7954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7956 = 9'hb0 == r_count_19_io_out ? io_r_176_b : _GEN_7955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7957 = 9'hb1 == r_count_19_io_out ? io_r_177_b : _GEN_7956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7958 = 9'hb2 == r_count_19_io_out ? io_r_178_b : _GEN_7957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7959 = 9'hb3 == r_count_19_io_out ? io_r_179_b : _GEN_7958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7960 = 9'hb4 == r_count_19_io_out ? io_r_180_b : _GEN_7959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7961 = 9'hb5 == r_count_19_io_out ? io_r_181_b : _GEN_7960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7962 = 9'hb6 == r_count_19_io_out ? io_r_182_b : _GEN_7961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7963 = 9'hb7 == r_count_19_io_out ? io_r_183_b : _GEN_7962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7964 = 9'hb8 == r_count_19_io_out ? io_r_184_b : _GEN_7963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7965 = 9'hb9 == r_count_19_io_out ? io_r_185_b : _GEN_7964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7966 = 9'hba == r_count_19_io_out ? io_r_186_b : _GEN_7965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7967 = 9'hbb == r_count_19_io_out ? io_r_187_b : _GEN_7966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7968 = 9'hbc == r_count_19_io_out ? io_r_188_b : _GEN_7967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7969 = 9'hbd == r_count_19_io_out ? io_r_189_b : _GEN_7968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7970 = 9'hbe == r_count_19_io_out ? io_r_190_b : _GEN_7969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7971 = 9'hbf == r_count_19_io_out ? io_r_191_b : _GEN_7970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7972 = 9'hc0 == r_count_19_io_out ? io_r_192_b : _GEN_7971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7973 = 9'hc1 == r_count_19_io_out ? io_r_193_b : _GEN_7972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7974 = 9'hc2 == r_count_19_io_out ? io_r_194_b : _GEN_7973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7975 = 9'hc3 == r_count_19_io_out ? io_r_195_b : _GEN_7974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7976 = 9'hc4 == r_count_19_io_out ? io_r_196_b : _GEN_7975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7977 = 9'hc5 == r_count_19_io_out ? io_r_197_b : _GEN_7976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7978 = 9'hc6 == r_count_19_io_out ? io_r_198_b : _GEN_7977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7979 = 9'hc7 == r_count_19_io_out ? io_r_199_b : _GEN_7978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7980 = 9'hc8 == r_count_19_io_out ? io_r_200_b : _GEN_7979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7981 = 9'hc9 == r_count_19_io_out ? io_r_201_b : _GEN_7980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7982 = 9'hca == r_count_19_io_out ? io_r_202_b : _GEN_7981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7983 = 9'hcb == r_count_19_io_out ? io_r_203_b : _GEN_7982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7984 = 9'hcc == r_count_19_io_out ? io_r_204_b : _GEN_7983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7985 = 9'hcd == r_count_19_io_out ? io_r_205_b : _GEN_7984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7986 = 9'hce == r_count_19_io_out ? io_r_206_b : _GEN_7985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7987 = 9'hcf == r_count_19_io_out ? io_r_207_b : _GEN_7986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7988 = 9'hd0 == r_count_19_io_out ? io_r_208_b : _GEN_7987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7989 = 9'hd1 == r_count_19_io_out ? io_r_209_b : _GEN_7988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7990 = 9'hd2 == r_count_19_io_out ? io_r_210_b : _GEN_7989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7991 = 9'hd3 == r_count_19_io_out ? io_r_211_b : _GEN_7990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7992 = 9'hd4 == r_count_19_io_out ? io_r_212_b : _GEN_7991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7993 = 9'hd5 == r_count_19_io_out ? io_r_213_b : _GEN_7992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7994 = 9'hd6 == r_count_19_io_out ? io_r_214_b : _GEN_7993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7995 = 9'hd7 == r_count_19_io_out ? io_r_215_b : _GEN_7994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7996 = 9'hd8 == r_count_19_io_out ? io_r_216_b : _GEN_7995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7997 = 9'hd9 == r_count_19_io_out ? io_r_217_b : _GEN_7996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7998 = 9'hda == r_count_19_io_out ? io_r_218_b : _GEN_7997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7999 = 9'hdb == r_count_19_io_out ? io_r_219_b : _GEN_7998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8000 = 9'hdc == r_count_19_io_out ? io_r_220_b : _GEN_7999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8001 = 9'hdd == r_count_19_io_out ? io_r_221_b : _GEN_8000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8002 = 9'hde == r_count_19_io_out ? io_r_222_b : _GEN_8001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8003 = 9'hdf == r_count_19_io_out ? io_r_223_b : _GEN_8002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8004 = 9'he0 == r_count_19_io_out ? io_r_224_b : _GEN_8003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8005 = 9'he1 == r_count_19_io_out ? io_r_225_b : _GEN_8004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8006 = 9'he2 == r_count_19_io_out ? io_r_226_b : _GEN_8005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8007 = 9'he3 == r_count_19_io_out ? io_r_227_b : _GEN_8006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8008 = 9'he4 == r_count_19_io_out ? io_r_228_b : _GEN_8007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8009 = 9'he5 == r_count_19_io_out ? io_r_229_b : _GEN_8008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8010 = 9'he6 == r_count_19_io_out ? io_r_230_b : _GEN_8009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8011 = 9'he7 == r_count_19_io_out ? io_r_231_b : _GEN_8010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8012 = 9'he8 == r_count_19_io_out ? io_r_232_b : _GEN_8011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8013 = 9'he9 == r_count_19_io_out ? io_r_233_b : _GEN_8012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8014 = 9'hea == r_count_19_io_out ? io_r_234_b : _GEN_8013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8015 = 9'heb == r_count_19_io_out ? io_r_235_b : _GEN_8014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8016 = 9'hec == r_count_19_io_out ? io_r_236_b : _GEN_8015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8017 = 9'hed == r_count_19_io_out ? io_r_237_b : _GEN_8016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8018 = 9'hee == r_count_19_io_out ? io_r_238_b : _GEN_8017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8019 = 9'hef == r_count_19_io_out ? io_r_239_b : _GEN_8018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8020 = 9'hf0 == r_count_19_io_out ? io_r_240_b : _GEN_8019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8021 = 9'hf1 == r_count_19_io_out ? io_r_241_b : _GEN_8020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8022 = 9'hf2 == r_count_19_io_out ? io_r_242_b : _GEN_8021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8023 = 9'hf3 == r_count_19_io_out ? io_r_243_b : _GEN_8022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8024 = 9'hf4 == r_count_19_io_out ? io_r_244_b : _GEN_8023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8025 = 9'hf5 == r_count_19_io_out ? io_r_245_b : _GEN_8024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8026 = 9'hf6 == r_count_19_io_out ? io_r_246_b : _GEN_8025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8027 = 9'hf7 == r_count_19_io_out ? io_r_247_b : _GEN_8026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8028 = 9'hf8 == r_count_19_io_out ? io_r_248_b : _GEN_8027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8029 = 9'hf9 == r_count_19_io_out ? io_r_249_b : _GEN_8028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8030 = 9'hfa == r_count_19_io_out ? io_r_250_b : _GEN_8029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8031 = 9'hfb == r_count_19_io_out ? io_r_251_b : _GEN_8030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8032 = 9'hfc == r_count_19_io_out ? io_r_252_b : _GEN_8031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8033 = 9'hfd == r_count_19_io_out ? io_r_253_b : _GEN_8032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8034 = 9'hfe == r_count_19_io_out ? io_r_254_b : _GEN_8033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8035 = 9'hff == r_count_19_io_out ? io_r_255_b : _GEN_8034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8036 = 9'h100 == r_count_19_io_out ? io_r_256_b : _GEN_8035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8037 = 9'h101 == r_count_19_io_out ? io_r_257_b : _GEN_8036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8038 = 9'h102 == r_count_19_io_out ? io_r_258_b : _GEN_8037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8039 = 9'h103 == r_count_19_io_out ? io_r_259_b : _GEN_8038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8040 = 9'h104 == r_count_19_io_out ? io_r_260_b : _GEN_8039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8041 = 9'h105 == r_count_19_io_out ? io_r_261_b : _GEN_8040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8042 = 9'h106 == r_count_19_io_out ? io_r_262_b : _GEN_8041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8043 = 9'h107 == r_count_19_io_out ? io_r_263_b : _GEN_8042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8044 = 9'h108 == r_count_19_io_out ? io_r_264_b : _GEN_8043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8045 = 9'h109 == r_count_19_io_out ? io_r_265_b : _GEN_8044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8046 = 9'h10a == r_count_19_io_out ? io_r_266_b : _GEN_8045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8047 = 9'h10b == r_count_19_io_out ? io_r_267_b : _GEN_8046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8048 = 9'h10c == r_count_19_io_out ? io_r_268_b : _GEN_8047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8049 = 9'h10d == r_count_19_io_out ? io_r_269_b : _GEN_8048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8050 = 9'h10e == r_count_19_io_out ? io_r_270_b : _GEN_8049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8051 = 9'h10f == r_count_19_io_out ? io_r_271_b : _GEN_8050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8052 = 9'h110 == r_count_19_io_out ? io_r_272_b : _GEN_8051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8053 = 9'h111 == r_count_19_io_out ? io_r_273_b : _GEN_8052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8054 = 9'h112 == r_count_19_io_out ? io_r_274_b : _GEN_8053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8055 = 9'h113 == r_count_19_io_out ? io_r_275_b : _GEN_8054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8056 = 9'h114 == r_count_19_io_out ? io_r_276_b : _GEN_8055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8057 = 9'h115 == r_count_19_io_out ? io_r_277_b : _GEN_8056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8058 = 9'h116 == r_count_19_io_out ? io_r_278_b : _GEN_8057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8059 = 9'h117 == r_count_19_io_out ? io_r_279_b : _GEN_8058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8060 = 9'h118 == r_count_19_io_out ? io_r_280_b : _GEN_8059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8061 = 9'h119 == r_count_19_io_out ? io_r_281_b : _GEN_8060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8062 = 9'h11a == r_count_19_io_out ? io_r_282_b : _GEN_8061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8063 = 9'h11b == r_count_19_io_out ? io_r_283_b : _GEN_8062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8064 = 9'h11c == r_count_19_io_out ? io_r_284_b : _GEN_8063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8065 = 9'h11d == r_count_19_io_out ? io_r_285_b : _GEN_8064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8066 = 9'h11e == r_count_19_io_out ? io_r_286_b : _GEN_8065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8067 = 9'h11f == r_count_19_io_out ? io_r_287_b : _GEN_8066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8068 = 9'h120 == r_count_19_io_out ? io_r_288_b : _GEN_8067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8069 = 9'h121 == r_count_19_io_out ? io_r_289_b : _GEN_8068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8070 = 9'h122 == r_count_19_io_out ? io_r_290_b : _GEN_8069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8071 = 9'h123 == r_count_19_io_out ? io_r_291_b : _GEN_8070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8072 = 9'h124 == r_count_19_io_out ? io_r_292_b : _GEN_8071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8073 = 9'h125 == r_count_19_io_out ? io_r_293_b : _GEN_8072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8074 = 9'h126 == r_count_19_io_out ? io_r_294_b : _GEN_8073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8075 = 9'h127 == r_count_19_io_out ? io_r_295_b : _GEN_8074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8076 = 9'h128 == r_count_19_io_out ? io_r_296_b : _GEN_8075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8077 = 9'h129 == r_count_19_io_out ? io_r_297_b : _GEN_8076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8078 = 9'h12a == r_count_19_io_out ? io_r_298_b : _GEN_8077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8079 = 9'h12b == r_count_19_io_out ? io_r_299_b : _GEN_8078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8080 = 9'h12c == r_count_19_io_out ? io_r_300_b : _GEN_8079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8081 = 9'h12d == r_count_19_io_out ? io_r_301_b : _GEN_8080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8082 = 9'h12e == r_count_19_io_out ? io_r_302_b : _GEN_8081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8083 = 9'h12f == r_count_19_io_out ? io_r_303_b : _GEN_8082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8084 = 9'h130 == r_count_19_io_out ? io_r_304_b : _GEN_8083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8085 = 9'h131 == r_count_19_io_out ? io_r_305_b : _GEN_8084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8086 = 9'h132 == r_count_19_io_out ? io_r_306_b : _GEN_8085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8087 = 9'h133 == r_count_19_io_out ? io_r_307_b : _GEN_8086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8088 = 9'h134 == r_count_19_io_out ? io_r_308_b : _GEN_8087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8089 = 9'h135 == r_count_19_io_out ? io_r_309_b : _GEN_8088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8090 = 9'h136 == r_count_19_io_out ? io_r_310_b : _GEN_8089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8091 = 9'h137 == r_count_19_io_out ? io_r_311_b : _GEN_8090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8092 = 9'h138 == r_count_19_io_out ? io_r_312_b : _GEN_8091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8093 = 9'h139 == r_count_19_io_out ? io_r_313_b : _GEN_8092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8094 = 9'h13a == r_count_19_io_out ? io_r_314_b : _GEN_8093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8095 = 9'h13b == r_count_19_io_out ? io_r_315_b : _GEN_8094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8096 = 9'h13c == r_count_19_io_out ? io_r_316_b : _GEN_8095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8097 = 9'h13d == r_count_19_io_out ? io_r_317_b : _GEN_8096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8098 = 9'h13e == r_count_19_io_out ? io_r_318_b : _GEN_8097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8099 = 9'h13f == r_count_19_io_out ? io_r_319_b : _GEN_8098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8100 = 9'h140 == r_count_19_io_out ? io_r_320_b : _GEN_8099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8101 = 9'h141 == r_count_19_io_out ? io_r_321_b : _GEN_8100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8102 = 9'h142 == r_count_19_io_out ? io_r_322_b : _GEN_8101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8103 = 9'h143 == r_count_19_io_out ? io_r_323_b : _GEN_8102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8104 = 9'h144 == r_count_19_io_out ? io_r_324_b : _GEN_8103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8105 = 9'h145 == r_count_19_io_out ? io_r_325_b : _GEN_8104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8106 = 9'h146 == r_count_19_io_out ? io_r_326_b : _GEN_8105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8107 = 9'h147 == r_count_19_io_out ? io_r_327_b : _GEN_8106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8108 = 9'h148 == r_count_19_io_out ? io_r_328_b : _GEN_8107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8109 = 9'h149 == r_count_19_io_out ? io_r_329_b : _GEN_8108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8110 = 9'h14a == r_count_19_io_out ? io_r_330_b : _GEN_8109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8111 = 9'h14b == r_count_19_io_out ? io_r_331_b : _GEN_8110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8112 = 9'h14c == r_count_19_io_out ? io_r_332_b : _GEN_8111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8113 = 9'h14d == r_count_19_io_out ? io_r_333_b : _GEN_8112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8114 = 9'h14e == r_count_19_io_out ? io_r_334_b : _GEN_8113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8115 = 9'h14f == r_count_19_io_out ? io_r_335_b : _GEN_8114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8116 = 9'h150 == r_count_19_io_out ? io_r_336_b : _GEN_8115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8117 = 9'h151 == r_count_19_io_out ? io_r_337_b : _GEN_8116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8118 = 9'h152 == r_count_19_io_out ? io_r_338_b : _GEN_8117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8119 = 9'h153 == r_count_19_io_out ? io_r_339_b : _GEN_8118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8120 = 9'h154 == r_count_19_io_out ? io_r_340_b : _GEN_8119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8121 = 9'h155 == r_count_19_io_out ? io_r_341_b : _GEN_8120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8122 = 9'h156 == r_count_19_io_out ? io_r_342_b : _GEN_8121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8123 = 9'h157 == r_count_19_io_out ? io_r_343_b : _GEN_8122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8124 = 9'h158 == r_count_19_io_out ? io_r_344_b : _GEN_8123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8125 = 9'h159 == r_count_19_io_out ? io_r_345_b : _GEN_8124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8126 = 9'h15a == r_count_19_io_out ? io_r_346_b : _GEN_8125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8127 = 9'h15b == r_count_19_io_out ? io_r_347_b : _GEN_8126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8128 = 9'h15c == r_count_19_io_out ? io_r_348_b : _GEN_8127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8129 = 9'h15d == r_count_19_io_out ? io_r_349_b : _GEN_8128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8130 = 9'h15e == r_count_19_io_out ? io_r_350_b : _GEN_8129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8131 = 9'h15f == r_count_19_io_out ? io_r_351_b : _GEN_8130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8132 = 9'h160 == r_count_19_io_out ? io_r_352_b : _GEN_8131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8133 = 9'h161 == r_count_19_io_out ? io_r_353_b : _GEN_8132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8134 = 9'h162 == r_count_19_io_out ? io_r_354_b : _GEN_8133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8135 = 9'h163 == r_count_19_io_out ? io_r_355_b : _GEN_8134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8136 = 9'h164 == r_count_19_io_out ? io_r_356_b : _GEN_8135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8137 = 9'h165 == r_count_19_io_out ? io_r_357_b : _GEN_8136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8138 = 9'h166 == r_count_19_io_out ? io_r_358_b : _GEN_8137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8139 = 9'h167 == r_count_19_io_out ? io_r_359_b : _GEN_8138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8140 = 9'h168 == r_count_19_io_out ? io_r_360_b : _GEN_8139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8141 = 9'h169 == r_count_19_io_out ? io_r_361_b : _GEN_8140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8142 = 9'h16a == r_count_19_io_out ? io_r_362_b : _GEN_8141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8143 = 9'h16b == r_count_19_io_out ? io_r_363_b : _GEN_8142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8144 = 9'h16c == r_count_19_io_out ? io_r_364_b : _GEN_8143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8145 = 9'h16d == r_count_19_io_out ? io_r_365_b : _GEN_8144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8146 = 9'h16e == r_count_19_io_out ? io_r_366_b : _GEN_8145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8147 = 9'h16f == r_count_19_io_out ? io_r_367_b : _GEN_8146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8148 = 9'h170 == r_count_19_io_out ? io_r_368_b : _GEN_8147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8149 = 9'h171 == r_count_19_io_out ? io_r_369_b : _GEN_8148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8150 = 9'h172 == r_count_19_io_out ? io_r_370_b : _GEN_8149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8151 = 9'h173 == r_count_19_io_out ? io_r_371_b : _GEN_8150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8152 = 9'h174 == r_count_19_io_out ? io_r_372_b : _GEN_8151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8153 = 9'h175 == r_count_19_io_out ? io_r_373_b : _GEN_8152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8154 = 9'h176 == r_count_19_io_out ? io_r_374_b : _GEN_8153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8155 = 9'h177 == r_count_19_io_out ? io_r_375_b : _GEN_8154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8156 = 9'h178 == r_count_19_io_out ? io_r_376_b : _GEN_8155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8157 = 9'h179 == r_count_19_io_out ? io_r_377_b : _GEN_8156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8158 = 9'h17a == r_count_19_io_out ? io_r_378_b : _GEN_8157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8159 = 9'h17b == r_count_19_io_out ? io_r_379_b : _GEN_8158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8160 = 9'h17c == r_count_19_io_out ? io_r_380_b : _GEN_8159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8161 = 9'h17d == r_count_19_io_out ? io_r_381_b : _GEN_8160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8162 = 9'h17e == r_count_19_io_out ? io_r_382_b : _GEN_8161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8163 = 9'h17f == r_count_19_io_out ? io_r_383_b : _GEN_8162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8164 = 9'h180 == r_count_19_io_out ? io_r_384_b : _GEN_8163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8165 = 9'h181 == r_count_19_io_out ? io_r_385_b : _GEN_8164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8166 = 9'h182 == r_count_19_io_out ? io_r_386_b : _GEN_8165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8167 = 9'h183 == r_count_19_io_out ? io_r_387_b : _GEN_8166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8168 = 9'h184 == r_count_19_io_out ? io_r_388_b : _GEN_8167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8169 = 9'h185 == r_count_19_io_out ? io_r_389_b : _GEN_8168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8170 = 9'h186 == r_count_19_io_out ? io_r_390_b : _GEN_8169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8171 = 9'h187 == r_count_19_io_out ? io_r_391_b : _GEN_8170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8172 = 9'h188 == r_count_19_io_out ? io_r_392_b : _GEN_8171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8173 = 9'h189 == r_count_19_io_out ? io_r_393_b : _GEN_8172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8174 = 9'h18a == r_count_19_io_out ? io_r_394_b : _GEN_8173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8175 = 9'h18b == r_count_19_io_out ? io_r_395_b : _GEN_8174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8176 = 9'h18c == r_count_19_io_out ? io_r_396_b : _GEN_8175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8177 = 9'h18d == r_count_19_io_out ? io_r_397_b : _GEN_8176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8178 = 9'h18e == r_count_19_io_out ? io_r_398_b : _GEN_8177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8181 = 9'h1 == r_count_20_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8182 = 9'h2 == r_count_20_io_out ? io_r_2_b : _GEN_8181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8183 = 9'h3 == r_count_20_io_out ? io_r_3_b : _GEN_8182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8184 = 9'h4 == r_count_20_io_out ? io_r_4_b : _GEN_8183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8185 = 9'h5 == r_count_20_io_out ? io_r_5_b : _GEN_8184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8186 = 9'h6 == r_count_20_io_out ? io_r_6_b : _GEN_8185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8187 = 9'h7 == r_count_20_io_out ? io_r_7_b : _GEN_8186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8188 = 9'h8 == r_count_20_io_out ? io_r_8_b : _GEN_8187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8189 = 9'h9 == r_count_20_io_out ? io_r_9_b : _GEN_8188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8190 = 9'ha == r_count_20_io_out ? io_r_10_b : _GEN_8189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8191 = 9'hb == r_count_20_io_out ? io_r_11_b : _GEN_8190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8192 = 9'hc == r_count_20_io_out ? io_r_12_b : _GEN_8191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8193 = 9'hd == r_count_20_io_out ? io_r_13_b : _GEN_8192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8194 = 9'he == r_count_20_io_out ? io_r_14_b : _GEN_8193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8195 = 9'hf == r_count_20_io_out ? io_r_15_b : _GEN_8194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8196 = 9'h10 == r_count_20_io_out ? io_r_16_b : _GEN_8195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8197 = 9'h11 == r_count_20_io_out ? io_r_17_b : _GEN_8196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8198 = 9'h12 == r_count_20_io_out ? io_r_18_b : _GEN_8197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8199 = 9'h13 == r_count_20_io_out ? io_r_19_b : _GEN_8198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8200 = 9'h14 == r_count_20_io_out ? io_r_20_b : _GEN_8199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8201 = 9'h15 == r_count_20_io_out ? io_r_21_b : _GEN_8200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8202 = 9'h16 == r_count_20_io_out ? io_r_22_b : _GEN_8201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8203 = 9'h17 == r_count_20_io_out ? io_r_23_b : _GEN_8202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8204 = 9'h18 == r_count_20_io_out ? io_r_24_b : _GEN_8203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8205 = 9'h19 == r_count_20_io_out ? io_r_25_b : _GEN_8204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8206 = 9'h1a == r_count_20_io_out ? io_r_26_b : _GEN_8205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8207 = 9'h1b == r_count_20_io_out ? io_r_27_b : _GEN_8206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8208 = 9'h1c == r_count_20_io_out ? io_r_28_b : _GEN_8207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8209 = 9'h1d == r_count_20_io_out ? io_r_29_b : _GEN_8208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8210 = 9'h1e == r_count_20_io_out ? io_r_30_b : _GEN_8209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8211 = 9'h1f == r_count_20_io_out ? io_r_31_b : _GEN_8210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8212 = 9'h20 == r_count_20_io_out ? io_r_32_b : _GEN_8211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8213 = 9'h21 == r_count_20_io_out ? io_r_33_b : _GEN_8212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8214 = 9'h22 == r_count_20_io_out ? io_r_34_b : _GEN_8213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8215 = 9'h23 == r_count_20_io_out ? io_r_35_b : _GEN_8214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8216 = 9'h24 == r_count_20_io_out ? io_r_36_b : _GEN_8215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8217 = 9'h25 == r_count_20_io_out ? io_r_37_b : _GEN_8216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8218 = 9'h26 == r_count_20_io_out ? io_r_38_b : _GEN_8217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8219 = 9'h27 == r_count_20_io_out ? io_r_39_b : _GEN_8218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8220 = 9'h28 == r_count_20_io_out ? io_r_40_b : _GEN_8219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8221 = 9'h29 == r_count_20_io_out ? io_r_41_b : _GEN_8220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8222 = 9'h2a == r_count_20_io_out ? io_r_42_b : _GEN_8221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8223 = 9'h2b == r_count_20_io_out ? io_r_43_b : _GEN_8222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8224 = 9'h2c == r_count_20_io_out ? io_r_44_b : _GEN_8223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8225 = 9'h2d == r_count_20_io_out ? io_r_45_b : _GEN_8224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8226 = 9'h2e == r_count_20_io_out ? io_r_46_b : _GEN_8225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8227 = 9'h2f == r_count_20_io_out ? io_r_47_b : _GEN_8226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8228 = 9'h30 == r_count_20_io_out ? io_r_48_b : _GEN_8227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8229 = 9'h31 == r_count_20_io_out ? io_r_49_b : _GEN_8228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8230 = 9'h32 == r_count_20_io_out ? io_r_50_b : _GEN_8229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8231 = 9'h33 == r_count_20_io_out ? io_r_51_b : _GEN_8230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8232 = 9'h34 == r_count_20_io_out ? io_r_52_b : _GEN_8231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8233 = 9'h35 == r_count_20_io_out ? io_r_53_b : _GEN_8232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8234 = 9'h36 == r_count_20_io_out ? io_r_54_b : _GEN_8233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8235 = 9'h37 == r_count_20_io_out ? io_r_55_b : _GEN_8234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8236 = 9'h38 == r_count_20_io_out ? io_r_56_b : _GEN_8235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8237 = 9'h39 == r_count_20_io_out ? io_r_57_b : _GEN_8236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8238 = 9'h3a == r_count_20_io_out ? io_r_58_b : _GEN_8237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8239 = 9'h3b == r_count_20_io_out ? io_r_59_b : _GEN_8238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8240 = 9'h3c == r_count_20_io_out ? io_r_60_b : _GEN_8239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8241 = 9'h3d == r_count_20_io_out ? io_r_61_b : _GEN_8240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8242 = 9'h3e == r_count_20_io_out ? io_r_62_b : _GEN_8241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8243 = 9'h3f == r_count_20_io_out ? io_r_63_b : _GEN_8242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8244 = 9'h40 == r_count_20_io_out ? io_r_64_b : _GEN_8243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8245 = 9'h41 == r_count_20_io_out ? io_r_65_b : _GEN_8244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8246 = 9'h42 == r_count_20_io_out ? io_r_66_b : _GEN_8245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8247 = 9'h43 == r_count_20_io_out ? io_r_67_b : _GEN_8246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8248 = 9'h44 == r_count_20_io_out ? io_r_68_b : _GEN_8247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8249 = 9'h45 == r_count_20_io_out ? io_r_69_b : _GEN_8248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8250 = 9'h46 == r_count_20_io_out ? io_r_70_b : _GEN_8249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8251 = 9'h47 == r_count_20_io_out ? io_r_71_b : _GEN_8250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8252 = 9'h48 == r_count_20_io_out ? io_r_72_b : _GEN_8251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8253 = 9'h49 == r_count_20_io_out ? io_r_73_b : _GEN_8252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8254 = 9'h4a == r_count_20_io_out ? io_r_74_b : _GEN_8253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8255 = 9'h4b == r_count_20_io_out ? io_r_75_b : _GEN_8254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8256 = 9'h4c == r_count_20_io_out ? io_r_76_b : _GEN_8255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8257 = 9'h4d == r_count_20_io_out ? io_r_77_b : _GEN_8256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8258 = 9'h4e == r_count_20_io_out ? io_r_78_b : _GEN_8257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8259 = 9'h4f == r_count_20_io_out ? io_r_79_b : _GEN_8258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8260 = 9'h50 == r_count_20_io_out ? io_r_80_b : _GEN_8259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8261 = 9'h51 == r_count_20_io_out ? io_r_81_b : _GEN_8260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8262 = 9'h52 == r_count_20_io_out ? io_r_82_b : _GEN_8261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8263 = 9'h53 == r_count_20_io_out ? io_r_83_b : _GEN_8262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8264 = 9'h54 == r_count_20_io_out ? io_r_84_b : _GEN_8263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8265 = 9'h55 == r_count_20_io_out ? io_r_85_b : _GEN_8264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8266 = 9'h56 == r_count_20_io_out ? io_r_86_b : _GEN_8265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8267 = 9'h57 == r_count_20_io_out ? io_r_87_b : _GEN_8266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8268 = 9'h58 == r_count_20_io_out ? io_r_88_b : _GEN_8267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8269 = 9'h59 == r_count_20_io_out ? io_r_89_b : _GEN_8268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8270 = 9'h5a == r_count_20_io_out ? io_r_90_b : _GEN_8269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8271 = 9'h5b == r_count_20_io_out ? io_r_91_b : _GEN_8270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8272 = 9'h5c == r_count_20_io_out ? io_r_92_b : _GEN_8271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8273 = 9'h5d == r_count_20_io_out ? io_r_93_b : _GEN_8272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8274 = 9'h5e == r_count_20_io_out ? io_r_94_b : _GEN_8273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8275 = 9'h5f == r_count_20_io_out ? io_r_95_b : _GEN_8274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8276 = 9'h60 == r_count_20_io_out ? io_r_96_b : _GEN_8275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8277 = 9'h61 == r_count_20_io_out ? io_r_97_b : _GEN_8276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8278 = 9'h62 == r_count_20_io_out ? io_r_98_b : _GEN_8277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8279 = 9'h63 == r_count_20_io_out ? io_r_99_b : _GEN_8278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8280 = 9'h64 == r_count_20_io_out ? io_r_100_b : _GEN_8279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8281 = 9'h65 == r_count_20_io_out ? io_r_101_b : _GEN_8280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8282 = 9'h66 == r_count_20_io_out ? io_r_102_b : _GEN_8281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8283 = 9'h67 == r_count_20_io_out ? io_r_103_b : _GEN_8282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8284 = 9'h68 == r_count_20_io_out ? io_r_104_b : _GEN_8283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8285 = 9'h69 == r_count_20_io_out ? io_r_105_b : _GEN_8284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8286 = 9'h6a == r_count_20_io_out ? io_r_106_b : _GEN_8285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8287 = 9'h6b == r_count_20_io_out ? io_r_107_b : _GEN_8286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8288 = 9'h6c == r_count_20_io_out ? io_r_108_b : _GEN_8287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8289 = 9'h6d == r_count_20_io_out ? io_r_109_b : _GEN_8288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8290 = 9'h6e == r_count_20_io_out ? io_r_110_b : _GEN_8289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8291 = 9'h6f == r_count_20_io_out ? io_r_111_b : _GEN_8290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8292 = 9'h70 == r_count_20_io_out ? io_r_112_b : _GEN_8291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8293 = 9'h71 == r_count_20_io_out ? io_r_113_b : _GEN_8292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8294 = 9'h72 == r_count_20_io_out ? io_r_114_b : _GEN_8293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8295 = 9'h73 == r_count_20_io_out ? io_r_115_b : _GEN_8294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8296 = 9'h74 == r_count_20_io_out ? io_r_116_b : _GEN_8295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8297 = 9'h75 == r_count_20_io_out ? io_r_117_b : _GEN_8296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8298 = 9'h76 == r_count_20_io_out ? io_r_118_b : _GEN_8297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8299 = 9'h77 == r_count_20_io_out ? io_r_119_b : _GEN_8298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8300 = 9'h78 == r_count_20_io_out ? io_r_120_b : _GEN_8299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8301 = 9'h79 == r_count_20_io_out ? io_r_121_b : _GEN_8300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8302 = 9'h7a == r_count_20_io_out ? io_r_122_b : _GEN_8301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8303 = 9'h7b == r_count_20_io_out ? io_r_123_b : _GEN_8302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8304 = 9'h7c == r_count_20_io_out ? io_r_124_b : _GEN_8303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8305 = 9'h7d == r_count_20_io_out ? io_r_125_b : _GEN_8304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8306 = 9'h7e == r_count_20_io_out ? io_r_126_b : _GEN_8305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8307 = 9'h7f == r_count_20_io_out ? io_r_127_b : _GEN_8306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8308 = 9'h80 == r_count_20_io_out ? io_r_128_b : _GEN_8307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8309 = 9'h81 == r_count_20_io_out ? io_r_129_b : _GEN_8308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8310 = 9'h82 == r_count_20_io_out ? io_r_130_b : _GEN_8309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8311 = 9'h83 == r_count_20_io_out ? io_r_131_b : _GEN_8310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8312 = 9'h84 == r_count_20_io_out ? io_r_132_b : _GEN_8311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8313 = 9'h85 == r_count_20_io_out ? io_r_133_b : _GEN_8312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8314 = 9'h86 == r_count_20_io_out ? io_r_134_b : _GEN_8313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8315 = 9'h87 == r_count_20_io_out ? io_r_135_b : _GEN_8314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8316 = 9'h88 == r_count_20_io_out ? io_r_136_b : _GEN_8315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8317 = 9'h89 == r_count_20_io_out ? io_r_137_b : _GEN_8316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8318 = 9'h8a == r_count_20_io_out ? io_r_138_b : _GEN_8317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8319 = 9'h8b == r_count_20_io_out ? io_r_139_b : _GEN_8318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8320 = 9'h8c == r_count_20_io_out ? io_r_140_b : _GEN_8319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8321 = 9'h8d == r_count_20_io_out ? io_r_141_b : _GEN_8320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8322 = 9'h8e == r_count_20_io_out ? io_r_142_b : _GEN_8321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8323 = 9'h8f == r_count_20_io_out ? io_r_143_b : _GEN_8322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8324 = 9'h90 == r_count_20_io_out ? io_r_144_b : _GEN_8323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8325 = 9'h91 == r_count_20_io_out ? io_r_145_b : _GEN_8324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8326 = 9'h92 == r_count_20_io_out ? io_r_146_b : _GEN_8325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8327 = 9'h93 == r_count_20_io_out ? io_r_147_b : _GEN_8326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8328 = 9'h94 == r_count_20_io_out ? io_r_148_b : _GEN_8327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8329 = 9'h95 == r_count_20_io_out ? io_r_149_b : _GEN_8328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8330 = 9'h96 == r_count_20_io_out ? io_r_150_b : _GEN_8329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8331 = 9'h97 == r_count_20_io_out ? io_r_151_b : _GEN_8330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8332 = 9'h98 == r_count_20_io_out ? io_r_152_b : _GEN_8331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8333 = 9'h99 == r_count_20_io_out ? io_r_153_b : _GEN_8332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8334 = 9'h9a == r_count_20_io_out ? io_r_154_b : _GEN_8333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8335 = 9'h9b == r_count_20_io_out ? io_r_155_b : _GEN_8334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8336 = 9'h9c == r_count_20_io_out ? io_r_156_b : _GEN_8335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8337 = 9'h9d == r_count_20_io_out ? io_r_157_b : _GEN_8336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8338 = 9'h9e == r_count_20_io_out ? io_r_158_b : _GEN_8337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8339 = 9'h9f == r_count_20_io_out ? io_r_159_b : _GEN_8338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8340 = 9'ha0 == r_count_20_io_out ? io_r_160_b : _GEN_8339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8341 = 9'ha1 == r_count_20_io_out ? io_r_161_b : _GEN_8340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8342 = 9'ha2 == r_count_20_io_out ? io_r_162_b : _GEN_8341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8343 = 9'ha3 == r_count_20_io_out ? io_r_163_b : _GEN_8342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8344 = 9'ha4 == r_count_20_io_out ? io_r_164_b : _GEN_8343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8345 = 9'ha5 == r_count_20_io_out ? io_r_165_b : _GEN_8344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8346 = 9'ha6 == r_count_20_io_out ? io_r_166_b : _GEN_8345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8347 = 9'ha7 == r_count_20_io_out ? io_r_167_b : _GEN_8346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8348 = 9'ha8 == r_count_20_io_out ? io_r_168_b : _GEN_8347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8349 = 9'ha9 == r_count_20_io_out ? io_r_169_b : _GEN_8348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8350 = 9'haa == r_count_20_io_out ? io_r_170_b : _GEN_8349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8351 = 9'hab == r_count_20_io_out ? io_r_171_b : _GEN_8350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8352 = 9'hac == r_count_20_io_out ? io_r_172_b : _GEN_8351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8353 = 9'had == r_count_20_io_out ? io_r_173_b : _GEN_8352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8354 = 9'hae == r_count_20_io_out ? io_r_174_b : _GEN_8353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8355 = 9'haf == r_count_20_io_out ? io_r_175_b : _GEN_8354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8356 = 9'hb0 == r_count_20_io_out ? io_r_176_b : _GEN_8355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8357 = 9'hb1 == r_count_20_io_out ? io_r_177_b : _GEN_8356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8358 = 9'hb2 == r_count_20_io_out ? io_r_178_b : _GEN_8357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8359 = 9'hb3 == r_count_20_io_out ? io_r_179_b : _GEN_8358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8360 = 9'hb4 == r_count_20_io_out ? io_r_180_b : _GEN_8359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8361 = 9'hb5 == r_count_20_io_out ? io_r_181_b : _GEN_8360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8362 = 9'hb6 == r_count_20_io_out ? io_r_182_b : _GEN_8361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8363 = 9'hb7 == r_count_20_io_out ? io_r_183_b : _GEN_8362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8364 = 9'hb8 == r_count_20_io_out ? io_r_184_b : _GEN_8363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8365 = 9'hb9 == r_count_20_io_out ? io_r_185_b : _GEN_8364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8366 = 9'hba == r_count_20_io_out ? io_r_186_b : _GEN_8365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8367 = 9'hbb == r_count_20_io_out ? io_r_187_b : _GEN_8366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8368 = 9'hbc == r_count_20_io_out ? io_r_188_b : _GEN_8367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8369 = 9'hbd == r_count_20_io_out ? io_r_189_b : _GEN_8368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8370 = 9'hbe == r_count_20_io_out ? io_r_190_b : _GEN_8369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8371 = 9'hbf == r_count_20_io_out ? io_r_191_b : _GEN_8370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8372 = 9'hc0 == r_count_20_io_out ? io_r_192_b : _GEN_8371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8373 = 9'hc1 == r_count_20_io_out ? io_r_193_b : _GEN_8372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8374 = 9'hc2 == r_count_20_io_out ? io_r_194_b : _GEN_8373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8375 = 9'hc3 == r_count_20_io_out ? io_r_195_b : _GEN_8374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8376 = 9'hc4 == r_count_20_io_out ? io_r_196_b : _GEN_8375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8377 = 9'hc5 == r_count_20_io_out ? io_r_197_b : _GEN_8376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8378 = 9'hc6 == r_count_20_io_out ? io_r_198_b : _GEN_8377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8379 = 9'hc7 == r_count_20_io_out ? io_r_199_b : _GEN_8378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8380 = 9'hc8 == r_count_20_io_out ? io_r_200_b : _GEN_8379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8381 = 9'hc9 == r_count_20_io_out ? io_r_201_b : _GEN_8380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8382 = 9'hca == r_count_20_io_out ? io_r_202_b : _GEN_8381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8383 = 9'hcb == r_count_20_io_out ? io_r_203_b : _GEN_8382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8384 = 9'hcc == r_count_20_io_out ? io_r_204_b : _GEN_8383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8385 = 9'hcd == r_count_20_io_out ? io_r_205_b : _GEN_8384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8386 = 9'hce == r_count_20_io_out ? io_r_206_b : _GEN_8385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8387 = 9'hcf == r_count_20_io_out ? io_r_207_b : _GEN_8386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8388 = 9'hd0 == r_count_20_io_out ? io_r_208_b : _GEN_8387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8389 = 9'hd1 == r_count_20_io_out ? io_r_209_b : _GEN_8388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8390 = 9'hd2 == r_count_20_io_out ? io_r_210_b : _GEN_8389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8391 = 9'hd3 == r_count_20_io_out ? io_r_211_b : _GEN_8390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8392 = 9'hd4 == r_count_20_io_out ? io_r_212_b : _GEN_8391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8393 = 9'hd5 == r_count_20_io_out ? io_r_213_b : _GEN_8392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8394 = 9'hd6 == r_count_20_io_out ? io_r_214_b : _GEN_8393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8395 = 9'hd7 == r_count_20_io_out ? io_r_215_b : _GEN_8394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8396 = 9'hd8 == r_count_20_io_out ? io_r_216_b : _GEN_8395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8397 = 9'hd9 == r_count_20_io_out ? io_r_217_b : _GEN_8396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8398 = 9'hda == r_count_20_io_out ? io_r_218_b : _GEN_8397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8399 = 9'hdb == r_count_20_io_out ? io_r_219_b : _GEN_8398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8400 = 9'hdc == r_count_20_io_out ? io_r_220_b : _GEN_8399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8401 = 9'hdd == r_count_20_io_out ? io_r_221_b : _GEN_8400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8402 = 9'hde == r_count_20_io_out ? io_r_222_b : _GEN_8401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8403 = 9'hdf == r_count_20_io_out ? io_r_223_b : _GEN_8402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8404 = 9'he0 == r_count_20_io_out ? io_r_224_b : _GEN_8403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8405 = 9'he1 == r_count_20_io_out ? io_r_225_b : _GEN_8404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8406 = 9'he2 == r_count_20_io_out ? io_r_226_b : _GEN_8405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8407 = 9'he3 == r_count_20_io_out ? io_r_227_b : _GEN_8406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8408 = 9'he4 == r_count_20_io_out ? io_r_228_b : _GEN_8407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8409 = 9'he5 == r_count_20_io_out ? io_r_229_b : _GEN_8408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8410 = 9'he6 == r_count_20_io_out ? io_r_230_b : _GEN_8409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8411 = 9'he7 == r_count_20_io_out ? io_r_231_b : _GEN_8410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8412 = 9'he8 == r_count_20_io_out ? io_r_232_b : _GEN_8411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8413 = 9'he9 == r_count_20_io_out ? io_r_233_b : _GEN_8412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8414 = 9'hea == r_count_20_io_out ? io_r_234_b : _GEN_8413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8415 = 9'heb == r_count_20_io_out ? io_r_235_b : _GEN_8414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8416 = 9'hec == r_count_20_io_out ? io_r_236_b : _GEN_8415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8417 = 9'hed == r_count_20_io_out ? io_r_237_b : _GEN_8416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8418 = 9'hee == r_count_20_io_out ? io_r_238_b : _GEN_8417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8419 = 9'hef == r_count_20_io_out ? io_r_239_b : _GEN_8418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8420 = 9'hf0 == r_count_20_io_out ? io_r_240_b : _GEN_8419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8421 = 9'hf1 == r_count_20_io_out ? io_r_241_b : _GEN_8420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8422 = 9'hf2 == r_count_20_io_out ? io_r_242_b : _GEN_8421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8423 = 9'hf3 == r_count_20_io_out ? io_r_243_b : _GEN_8422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8424 = 9'hf4 == r_count_20_io_out ? io_r_244_b : _GEN_8423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8425 = 9'hf5 == r_count_20_io_out ? io_r_245_b : _GEN_8424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8426 = 9'hf6 == r_count_20_io_out ? io_r_246_b : _GEN_8425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8427 = 9'hf7 == r_count_20_io_out ? io_r_247_b : _GEN_8426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8428 = 9'hf8 == r_count_20_io_out ? io_r_248_b : _GEN_8427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8429 = 9'hf9 == r_count_20_io_out ? io_r_249_b : _GEN_8428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8430 = 9'hfa == r_count_20_io_out ? io_r_250_b : _GEN_8429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8431 = 9'hfb == r_count_20_io_out ? io_r_251_b : _GEN_8430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8432 = 9'hfc == r_count_20_io_out ? io_r_252_b : _GEN_8431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8433 = 9'hfd == r_count_20_io_out ? io_r_253_b : _GEN_8432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8434 = 9'hfe == r_count_20_io_out ? io_r_254_b : _GEN_8433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8435 = 9'hff == r_count_20_io_out ? io_r_255_b : _GEN_8434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8436 = 9'h100 == r_count_20_io_out ? io_r_256_b : _GEN_8435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8437 = 9'h101 == r_count_20_io_out ? io_r_257_b : _GEN_8436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8438 = 9'h102 == r_count_20_io_out ? io_r_258_b : _GEN_8437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8439 = 9'h103 == r_count_20_io_out ? io_r_259_b : _GEN_8438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8440 = 9'h104 == r_count_20_io_out ? io_r_260_b : _GEN_8439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8441 = 9'h105 == r_count_20_io_out ? io_r_261_b : _GEN_8440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8442 = 9'h106 == r_count_20_io_out ? io_r_262_b : _GEN_8441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8443 = 9'h107 == r_count_20_io_out ? io_r_263_b : _GEN_8442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8444 = 9'h108 == r_count_20_io_out ? io_r_264_b : _GEN_8443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8445 = 9'h109 == r_count_20_io_out ? io_r_265_b : _GEN_8444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8446 = 9'h10a == r_count_20_io_out ? io_r_266_b : _GEN_8445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8447 = 9'h10b == r_count_20_io_out ? io_r_267_b : _GEN_8446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8448 = 9'h10c == r_count_20_io_out ? io_r_268_b : _GEN_8447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8449 = 9'h10d == r_count_20_io_out ? io_r_269_b : _GEN_8448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8450 = 9'h10e == r_count_20_io_out ? io_r_270_b : _GEN_8449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8451 = 9'h10f == r_count_20_io_out ? io_r_271_b : _GEN_8450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8452 = 9'h110 == r_count_20_io_out ? io_r_272_b : _GEN_8451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8453 = 9'h111 == r_count_20_io_out ? io_r_273_b : _GEN_8452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8454 = 9'h112 == r_count_20_io_out ? io_r_274_b : _GEN_8453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8455 = 9'h113 == r_count_20_io_out ? io_r_275_b : _GEN_8454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8456 = 9'h114 == r_count_20_io_out ? io_r_276_b : _GEN_8455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8457 = 9'h115 == r_count_20_io_out ? io_r_277_b : _GEN_8456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8458 = 9'h116 == r_count_20_io_out ? io_r_278_b : _GEN_8457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8459 = 9'h117 == r_count_20_io_out ? io_r_279_b : _GEN_8458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8460 = 9'h118 == r_count_20_io_out ? io_r_280_b : _GEN_8459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8461 = 9'h119 == r_count_20_io_out ? io_r_281_b : _GEN_8460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8462 = 9'h11a == r_count_20_io_out ? io_r_282_b : _GEN_8461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8463 = 9'h11b == r_count_20_io_out ? io_r_283_b : _GEN_8462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8464 = 9'h11c == r_count_20_io_out ? io_r_284_b : _GEN_8463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8465 = 9'h11d == r_count_20_io_out ? io_r_285_b : _GEN_8464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8466 = 9'h11e == r_count_20_io_out ? io_r_286_b : _GEN_8465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8467 = 9'h11f == r_count_20_io_out ? io_r_287_b : _GEN_8466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8468 = 9'h120 == r_count_20_io_out ? io_r_288_b : _GEN_8467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8469 = 9'h121 == r_count_20_io_out ? io_r_289_b : _GEN_8468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8470 = 9'h122 == r_count_20_io_out ? io_r_290_b : _GEN_8469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8471 = 9'h123 == r_count_20_io_out ? io_r_291_b : _GEN_8470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8472 = 9'h124 == r_count_20_io_out ? io_r_292_b : _GEN_8471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8473 = 9'h125 == r_count_20_io_out ? io_r_293_b : _GEN_8472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8474 = 9'h126 == r_count_20_io_out ? io_r_294_b : _GEN_8473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8475 = 9'h127 == r_count_20_io_out ? io_r_295_b : _GEN_8474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8476 = 9'h128 == r_count_20_io_out ? io_r_296_b : _GEN_8475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8477 = 9'h129 == r_count_20_io_out ? io_r_297_b : _GEN_8476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8478 = 9'h12a == r_count_20_io_out ? io_r_298_b : _GEN_8477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8479 = 9'h12b == r_count_20_io_out ? io_r_299_b : _GEN_8478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8480 = 9'h12c == r_count_20_io_out ? io_r_300_b : _GEN_8479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8481 = 9'h12d == r_count_20_io_out ? io_r_301_b : _GEN_8480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8482 = 9'h12e == r_count_20_io_out ? io_r_302_b : _GEN_8481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8483 = 9'h12f == r_count_20_io_out ? io_r_303_b : _GEN_8482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8484 = 9'h130 == r_count_20_io_out ? io_r_304_b : _GEN_8483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8485 = 9'h131 == r_count_20_io_out ? io_r_305_b : _GEN_8484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8486 = 9'h132 == r_count_20_io_out ? io_r_306_b : _GEN_8485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8487 = 9'h133 == r_count_20_io_out ? io_r_307_b : _GEN_8486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8488 = 9'h134 == r_count_20_io_out ? io_r_308_b : _GEN_8487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8489 = 9'h135 == r_count_20_io_out ? io_r_309_b : _GEN_8488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8490 = 9'h136 == r_count_20_io_out ? io_r_310_b : _GEN_8489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8491 = 9'h137 == r_count_20_io_out ? io_r_311_b : _GEN_8490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8492 = 9'h138 == r_count_20_io_out ? io_r_312_b : _GEN_8491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8493 = 9'h139 == r_count_20_io_out ? io_r_313_b : _GEN_8492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8494 = 9'h13a == r_count_20_io_out ? io_r_314_b : _GEN_8493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8495 = 9'h13b == r_count_20_io_out ? io_r_315_b : _GEN_8494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8496 = 9'h13c == r_count_20_io_out ? io_r_316_b : _GEN_8495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8497 = 9'h13d == r_count_20_io_out ? io_r_317_b : _GEN_8496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8498 = 9'h13e == r_count_20_io_out ? io_r_318_b : _GEN_8497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8499 = 9'h13f == r_count_20_io_out ? io_r_319_b : _GEN_8498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8500 = 9'h140 == r_count_20_io_out ? io_r_320_b : _GEN_8499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8501 = 9'h141 == r_count_20_io_out ? io_r_321_b : _GEN_8500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8502 = 9'h142 == r_count_20_io_out ? io_r_322_b : _GEN_8501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8503 = 9'h143 == r_count_20_io_out ? io_r_323_b : _GEN_8502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8504 = 9'h144 == r_count_20_io_out ? io_r_324_b : _GEN_8503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8505 = 9'h145 == r_count_20_io_out ? io_r_325_b : _GEN_8504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8506 = 9'h146 == r_count_20_io_out ? io_r_326_b : _GEN_8505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8507 = 9'h147 == r_count_20_io_out ? io_r_327_b : _GEN_8506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8508 = 9'h148 == r_count_20_io_out ? io_r_328_b : _GEN_8507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8509 = 9'h149 == r_count_20_io_out ? io_r_329_b : _GEN_8508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8510 = 9'h14a == r_count_20_io_out ? io_r_330_b : _GEN_8509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8511 = 9'h14b == r_count_20_io_out ? io_r_331_b : _GEN_8510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8512 = 9'h14c == r_count_20_io_out ? io_r_332_b : _GEN_8511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8513 = 9'h14d == r_count_20_io_out ? io_r_333_b : _GEN_8512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8514 = 9'h14e == r_count_20_io_out ? io_r_334_b : _GEN_8513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8515 = 9'h14f == r_count_20_io_out ? io_r_335_b : _GEN_8514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8516 = 9'h150 == r_count_20_io_out ? io_r_336_b : _GEN_8515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8517 = 9'h151 == r_count_20_io_out ? io_r_337_b : _GEN_8516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8518 = 9'h152 == r_count_20_io_out ? io_r_338_b : _GEN_8517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8519 = 9'h153 == r_count_20_io_out ? io_r_339_b : _GEN_8518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8520 = 9'h154 == r_count_20_io_out ? io_r_340_b : _GEN_8519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8521 = 9'h155 == r_count_20_io_out ? io_r_341_b : _GEN_8520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8522 = 9'h156 == r_count_20_io_out ? io_r_342_b : _GEN_8521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8523 = 9'h157 == r_count_20_io_out ? io_r_343_b : _GEN_8522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8524 = 9'h158 == r_count_20_io_out ? io_r_344_b : _GEN_8523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8525 = 9'h159 == r_count_20_io_out ? io_r_345_b : _GEN_8524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8526 = 9'h15a == r_count_20_io_out ? io_r_346_b : _GEN_8525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8527 = 9'h15b == r_count_20_io_out ? io_r_347_b : _GEN_8526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8528 = 9'h15c == r_count_20_io_out ? io_r_348_b : _GEN_8527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8529 = 9'h15d == r_count_20_io_out ? io_r_349_b : _GEN_8528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8530 = 9'h15e == r_count_20_io_out ? io_r_350_b : _GEN_8529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8531 = 9'h15f == r_count_20_io_out ? io_r_351_b : _GEN_8530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8532 = 9'h160 == r_count_20_io_out ? io_r_352_b : _GEN_8531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8533 = 9'h161 == r_count_20_io_out ? io_r_353_b : _GEN_8532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8534 = 9'h162 == r_count_20_io_out ? io_r_354_b : _GEN_8533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8535 = 9'h163 == r_count_20_io_out ? io_r_355_b : _GEN_8534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8536 = 9'h164 == r_count_20_io_out ? io_r_356_b : _GEN_8535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8537 = 9'h165 == r_count_20_io_out ? io_r_357_b : _GEN_8536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8538 = 9'h166 == r_count_20_io_out ? io_r_358_b : _GEN_8537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8539 = 9'h167 == r_count_20_io_out ? io_r_359_b : _GEN_8538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8540 = 9'h168 == r_count_20_io_out ? io_r_360_b : _GEN_8539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8541 = 9'h169 == r_count_20_io_out ? io_r_361_b : _GEN_8540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8542 = 9'h16a == r_count_20_io_out ? io_r_362_b : _GEN_8541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8543 = 9'h16b == r_count_20_io_out ? io_r_363_b : _GEN_8542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8544 = 9'h16c == r_count_20_io_out ? io_r_364_b : _GEN_8543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8545 = 9'h16d == r_count_20_io_out ? io_r_365_b : _GEN_8544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8546 = 9'h16e == r_count_20_io_out ? io_r_366_b : _GEN_8545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8547 = 9'h16f == r_count_20_io_out ? io_r_367_b : _GEN_8546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8548 = 9'h170 == r_count_20_io_out ? io_r_368_b : _GEN_8547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8549 = 9'h171 == r_count_20_io_out ? io_r_369_b : _GEN_8548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8550 = 9'h172 == r_count_20_io_out ? io_r_370_b : _GEN_8549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8551 = 9'h173 == r_count_20_io_out ? io_r_371_b : _GEN_8550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8552 = 9'h174 == r_count_20_io_out ? io_r_372_b : _GEN_8551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8553 = 9'h175 == r_count_20_io_out ? io_r_373_b : _GEN_8552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8554 = 9'h176 == r_count_20_io_out ? io_r_374_b : _GEN_8553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8555 = 9'h177 == r_count_20_io_out ? io_r_375_b : _GEN_8554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8556 = 9'h178 == r_count_20_io_out ? io_r_376_b : _GEN_8555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8557 = 9'h179 == r_count_20_io_out ? io_r_377_b : _GEN_8556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8558 = 9'h17a == r_count_20_io_out ? io_r_378_b : _GEN_8557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8559 = 9'h17b == r_count_20_io_out ? io_r_379_b : _GEN_8558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8560 = 9'h17c == r_count_20_io_out ? io_r_380_b : _GEN_8559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8561 = 9'h17d == r_count_20_io_out ? io_r_381_b : _GEN_8560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8562 = 9'h17e == r_count_20_io_out ? io_r_382_b : _GEN_8561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8563 = 9'h17f == r_count_20_io_out ? io_r_383_b : _GEN_8562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8564 = 9'h180 == r_count_20_io_out ? io_r_384_b : _GEN_8563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8565 = 9'h181 == r_count_20_io_out ? io_r_385_b : _GEN_8564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8566 = 9'h182 == r_count_20_io_out ? io_r_386_b : _GEN_8565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8567 = 9'h183 == r_count_20_io_out ? io_r_387_b : _GEN_8566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8568 = 9'h184 == r_count_20_io_out ? io_r_388_b : _GEN_8567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8569 = 9'h185 == r_count_20_io_out ? io_r_389_b : _GEN_8568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8570 = 9'h186 == r_count_20_io_out ? io_r_390_b : _GEN_8569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8571 = 9'h187 == r_count_20_io_out ? io_r_391_b : _GEN_8570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8572 = 9'h188 == r_count_20_io_out ? io_r_392_b : _GEN_8571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8573 = 9'h189 == r_count_20_io_out ? io_r_393_b : _GEN_8572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8574 = 9'h18a == r_count_20_io_out ? io_r_394_b : _GEN_8573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8575 = 9'h18b == r_count_20_io_out ? io_r_395_b : _GEN_8574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8576 = 9'h18c == r_count_20_io_out ? io_r_396_b : _GEN_8575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8577 = 9'h18d == r_count_20_io_out ? io_r_397_b : _GEN_8576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8578 = 9'h18e == r_count_20_io_out ? io_r_398_b : _GEN_8577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8581 = 9'h1 == r_count_21_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8582 = 9'h2 == r_count_21_io_out ? io_r_2_b : _GEN_8581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8583 = 9'h3 == r_count_21_io_out ? io_r_3_b : _GEN_8582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8584 = 9'h4 == r_count_21_io_out ? io_r_4_b : _GEN_8583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8585 = 9'h5 == r_count_21_io_out ? io_r_5_b : _GEN_8584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8586 = 9'h6 == r_count_21_io_out ? io_r_6_b : _GEN_8585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8587 = 9'h7 == r_count_21_io_out ? io_r_7_b : _GEN_8586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8588 = 9'h8 == r_count_21_io_out ? io_r_8_b : _GEN_8587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8589 = 9'h9 == r_count_21_io_out ? io_r_9_b : _GEN_8588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8590 = 9'ha == r_count_21_io_out ? io_r_10_b : _GEN_8589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8591 = 9'hb == r_count_21_io_out ? io_r_11_b : _GEN_8590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8592 = 9'hc == r_count_21_io_out ? io_r_12_b : _GEN_8591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8593 = 9'hd == r_count_21_io_out ? io_r_13_b : _GEN_8592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8594 = 9'he == r_count_21_io_out ? io_r_14_b : _GEN_8593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8595 = 9'hf == r_count_21_io_out ? io_r_15_b : _GEN_8594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8596 = 9'h10 == r_count_21_io_out ? io_r_16_b : _GEN_8595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8597 = 9'h11 == r_count_21_io_out ? io_r_17_b : _GEN_8596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8598 = 9'h12 == r_count_21_io_out ? io_r_18_b : _GEN_8597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8599 = 9'h13 == r_count_21_io_out ? io_r_19_b : _GEN_8598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8600 = 9'h14 == r_count_21_io_out ? io_r_20_b : _GEN_8599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8601 = 9'h15 == r_count_21_io_out ? io_r_21_b : _GEN_8600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8602 = 9'h16 == r_count_21_io_out ? io_r_22_b : _GEN_8601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8603 = 9'h17 == r_count_21_io_out ? io_r_23_b : _GEN_8602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8604 = 9'h18 == r_count_21_io_out ? io_r_24_b : _GEN_8603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8605 = 9'h19 == r_count_21_io_out ? io_r_25_b : _GEN_8604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8606 = 9'h1a == r_count_21_io_out ? io_r_26_b : _GEN_8605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8607 = 9'h1b == r_count_21_io_out ? io_r_27_b : _GEN_8606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8608 = 9'h1c == r_count_21_io_out ? io_r_28_b : _GEN_8607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8609 = 9'h1d == r_count_21_io_out ? io_r_29_b : _GEN_8608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8610 = 9'h1e == r_count_21_io_out ? io_r_30_b : _GEN_8609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8611 = 9'h1f == r_count_21_io_out ? io_r_31_b : _GEN_8610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8612 = 9'h20 == r_count_21_io_out ? io_r_32_b : _GEN_8611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8613 = 9'h21 == r_count_21_io_out ? io_r_33_b : _GEN_8612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8614 = 9'h22 == r_count_21_io_out ? io_r_34_b : _GEN_8613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8615 = 9'h23 == r_count_21_io_out ? io_r_35_b : _GEN_8614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8616 = 9'h24 == r_count_21_io_out ? io_r_36_b : _GEN_8615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8617 = 9'h25 == r_count_21_io_out ? io_r_37_b : _GEN_8616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8618 = 9'h26 == r_count_21_io_out ? io_r_38_b : _GEN_8617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8619 = 9'h27 == r_count_21_io_out ? io_r_39_b : _GEN_8618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8620 = 9'h28 == r_count_21_io_out ? io_r_40_b : _GEN_8619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8621 = 9'h29 == r_count_21_io_out ? io_r_41_b : _GEN_8620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8622 = 9'h2a == r_count_21_io_out ? io_r_42_b : _GEN_8621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8623 = 9'h2b == r_count_21_io_out ? io_r_43_b : _GEN_8622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8624 = 9'h2c == r_count_21_io_out ? io_r_44_b : _GEN_8623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8625 = 9'h2d == r_count_21_io_out ? io_r_45_b : _GEN_8624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8626 = 9'h2e == r_count_21_io_out ? io_r_46_b : _GEN_8625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8627 = 9'h2f == r_count_21_io_out ? io_r_47_b : _GEN_8626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8628 = 9'h30 == r_count_21_io_out ? io_r_48_b : _GEN_8627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8629 = 9'h31 == r_count_21_io_out ? io_r_49_b : _GEN_8628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8630 = 9'h32 == r_count_21_io_out ? io_r_50_b : _GEN_8629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8631 = 9'h33 == r_count_21_io_out ? io_r_51_b : _GEN_8630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8632 = 9'h34 == r_count_21_io_out ? io_r_52_b : _GEN_8631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8633 = 9'h35 == r_count_21_io_out ? io_r_53_b : _GEN_8632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8634 = 9'h36 == r_count_21_io_out ? io_r_54_b : _GEN_8633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8635 = 9'h37 == r_count_21_io_out ? io_r_55_b : _GEN_8634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8636 = 9'h38 == r_count_21_io_out ? io_r_56_b : _GEN_8635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8637 = 9'h39 == r_count_21_io_out ? io_r_57_b : _GEN_8636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8638 = 9'h3a == r_count_21_io_out ? io_r_58_b : _GEN_8637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8639 = 9'h3b == r_count_21_io_out ? io_r_59_b : _GEN_8638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8640 = 9'h3c == r_count_21_io_out ? io_r_60_b : _GEN_8639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8641 = 9'h3d == r_count_21_io_out ? io_r_61_b : _GEN_8640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8642 = 9'h3e == r_count_21_io_out ? io_r_62_b : _GEN_8641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8643 = 9'h3f == r_count_21_io_out ? io_r_63_b : _GEN_8642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8644 = 9'h40 == r_count_21_io_out ? io_r_64_b : _GEN_8643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8645 = 9'h41 == r_count_21_io_out ? io_r_65_b : _GEN_8644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8646 = 9'h42 == r_count_21_io_out ? io_r_66_b : _GEN_8645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8647 = 9'h43 == r_count_21_io_out ? io_r_67_b : _GEN_8646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8648 = 9'h44 == r_count_21_io_out ? io_r_68_b : _GEN_8647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8649 = 9'h45 == r_count_21_io_out ? io_r_69_b : _GEN_8648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8650 = 9'h46 == r_count_21_io_out ? io_r_70_b : _GEN_8649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8651 = 9'h47 == r_count_21_io_out ? io_r_71_b : _GEN_8650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8652 = 9'h48 == r_count_21_io_out ? io_r_72_b : _GEN_8651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8653 = 9'h49 == r_count_21_io_out ? io_r_73_b : _GEN_8652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8654 = 9'h4a == r_count_21_io_out ? io_r_74_b : _GEN_8653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8655 = 9'h4b == r_count_21_io_out ? io_r_75_b : _GEN_8654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8656 = 9'h4c == r_count_21_io_out ? io_r_76_b : _GEN_8655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8657 = 9'h4d == r_count_21_io_out ? io_r_77_b : _GEN_8656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8658 = 9'h4e == r_count_21_io_out ? io_r_78_b : _GEN_8657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8659 = 9'h4f == r_count_21_io_out ? io_r_79_b : _GEN_8658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8660 = 9'h50 == r_count_21_io_out ? io_r_80_b : _GEN_8659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8661 = 9'h51 == r_count_21_io_out ? io_r_81_b : _GEN_8660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8662 = 9'h52 == r_count_21_io_out ? io_r_82_b : _GEN_8661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8663 = 9'h53 == r_count_21_io_out ? io_r_83_b : _GEN_8662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8664 = 9'h54 == r_count_21_io_out ? io_r_84_b : _GEN_8663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8665 = 9'h55 == r_count_21_io_out ? io_r_85_b : _GEN_8664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8666 = 9'h56 == r_count_21_io_out ? io_r_86_b : _GEN_8665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8667 = 9'h57 == r_count_21_io_out ? io_r_87_b : _GEN_8666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8668 = 9'h58 == r_count_21_io_out ? io_r_88_b : _GEN_8667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8669 = 9'h59 == r_count_21_io_out ? io_r_89_b : _GEN_8668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8670 = 9'h5a == r_count_21_io_out ? io_r_90_b : _GEN_8669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8671 = 9'h5b == r_count_21_io_out ? io_r_91_b : _GEN_8670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8672 = 9'h5c == r_count_21_io_out ? io_r_92_b : _GEN_8671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8673 = 9'h5d == r_count_21_io_out ? io_r_93_b : _GEN_8672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8674 = 9'h5e == r_count_21_io_out ? io_r_94_b : _GEN_8673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8675 = 9'h5f == r_count_21_io_out ? io_r_95_b : _GEN_8674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8676 = 9'h60 == r_count_21_io_out ? io_r_96_b : _GEN_8675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8677 = 9'h61 == r_count_21_io_out ? io_r_97_b : _GEN_8676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8678 = 9'h62 == r_count_21_io_out ? io_r_98_b : _GEN_8677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8679 = 9'h63 == r_count_21_io_out ? io_r_99_b : _GEN_8678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8680 = 9'h64 == r_count_21_io_out ? io_r_100_b : _GEN_8679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8681 = 9'h65 == r_count_21_io_out ? io_r_101_b : _GEN_8680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8682 = 9'h66 == r_count_21_io_out ? io_r_102_b : _GEN_8681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8683 = 9'h67 == r_count_21_io_out ? io_r_103_b : _GEN_8682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8684 = 9'h68 == r_count_21_io_out ? io_r_104_b : _GEN_8683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8685 = 9'h69 == r_count_21_io_out ? io_r_105_b : _GEN_8684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8686 = 9'h6a == r_count_21_io_out ? io_r_106_b : _GEN_8685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8687 = 9'h6b == r_count_21_io_out ? io_r_107_b : _GEN_8686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8688 = 9'h6c == r_count_21_io_out ? io_r_108_b : _GEN_8687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8689 = 9'h6d == r_count_21_io_out ? io_r_109_b : _GEN_8688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8690 = 9'h6e == r_count_21_io_out ? io_r_110_b : _GEN_8689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8691 = 9'h6f == r_count_21_io_out ? io_r_111_b : _GEN_8690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8692 = 9'h70 == r_count_21_io_out ? io_r_112_b : _GEN_8691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8693 = 9'h71 == r_count_21_io_out ? io_r_113_b : _GEN_8692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8694 = 9'h72 == r_count_21_io_out ? io_r_114_b : _GEN_8693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8695 = 9'h73 == r_count_21_io_out ? io_r_115_b : _GEN_8694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8696 = 9'h74 == r_count_21_io_out ? io_r_116_b : _GEN_8695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8697 = 9'h75 == r_count_21_io_out ? io_r_117_b : _GEN_8696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8698 = 9'h76 == r_count_21_io_out ? io_r_118_b : _GEN_8697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8699 = 9'h77 == r_count_21_io_out ? io_r_119_b : _GEN_8698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8700 = 9'h78 == r_count_21_io_out ? io_r_120_b : _GEN_8699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8701 = 9'h79 == r_count_21_io_out ? io_r_121_b : _GEN_8700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8702 = 9'h7a == r_count_21_io_out ? io_r_122_b : _GEN_8701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8703 = 9'h7b == r_count_21_io_out ? io_r_123_b : _GEN_8702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8704 = 9'h7c == r_count_21_io_out ? io_r_124_b : _GEN_8703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8705 = 9'h7d == r_count_21_io_out ? io_r_125_b : _GEN_8704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8706 = 9'h7e == r_count_21_io_out ? io_r_126_b : _GEN_8705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8707 = 9'h7f == r_count_21_io_out ? io_r_127_b : _GEN_8706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8708 = 9'h80 == r_count_21_io_out ? io_r_128_b : _GEN_8707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8709 = 9'h81 == r_count_21_io_out ? io_r_129_b : _GEN_8708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8710 = 9'h82 == r_count_21_io_out ? io_r_130_b : _GEN_8709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8711 = 9'h83 == r_count_21_io_out ? io_r_131_b : _GEN_8710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8712 = 9'h84 == r_count_21_io_out ? io_r_132_b : _GEN_8711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8713 = 9'h85 == r_count_21_io_out ? io_r_133_b : _GEN_8712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8714 = 9'h86 == r_count_21_io_out ? io_r_134_b : _GEN_8713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8715 = 9'h87 == r_count_21_io_out ? io_r_135_b : _GEN_8714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8716 = 9'h88 == r_count_21_io_out ? io_r_136_b : _GEN_8715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8717 = 9'h89 == r_count_21_io_out ? io_r_137_b : _GEN_8716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8718 = 9'h8a == r_count_21_io_out ? io_r_138_b : _GEN_8717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8719 = 9'h8b == r_count_21_io_out ? io_r_139_b : _GEN_8718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8720 = 9'h8c == r_count_21_io_out ? io_r_140_b : _GEN_8719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8721 = 9'h8d == r_count_21_io_out ? io_r_141_b : _GEN_8720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8722 = 9'h8e == r_count_21_io_out ? io_r_142_b : _GEN_8721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8723 = 9'h8f == r_count_21_io_out ? io_r_143_b : _GEN_8722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8724 = 9'h90 == r_count_21_io_out ? io_r_144_b : _GEN_8723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8725 = 9'h91 == r_count_21_io_out ? io_r_145_b : _GEN_8724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8726 = 9'h92 == r_count_21_io_out ? io_r_146_b : _GEN_8725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8727 = 9'h93 == r_count_21_io_out ? io_r_147_b : _GEN_8726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8728 = 9'h94 == r_count_21_io_out ? io_r_148_b : _GEN_8727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8729 = 9'h95 == r_count_21_io_out ? io_r_149_b : _GEN_8728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8730 = 9'h96 == r_count_21_io_out ? io_r_150_b : _GEN_8729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8731 = 9'h97 == r_count_21_io_out ? io_r_151_b : _GEN_8730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8732 = 9'h98 == r_count_21_io_out ? io_r_152_b : _GEN_8731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8733 = 9'h99 == r_count_21_io_out ? io_r_153_b : _GEN_8732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8734 = 9'h9a == r_count_21_io_out ? io_r_154_b : _GEN_8733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8735 = 9'h9b == r_count_21_io_out ? io_r_155_b : _GEN_8734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8736 = 9'h9c == r_count_21_io_out ? io_r_156_b : _GEN_8735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8737 = 9'h9d == r_count_21_io_out ? io_r_157_b : _GEN_8736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8738 = 9'h9e == r_count_21_io_out ? io_r_158_b : _GEN_8737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8739 = 9'h9f == r_count_21_io_out ? io_r_159_b : _GEN_8738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8740 = 9'ha0 == r_count_21_io_out ? io_r_160_b : _GEN_8739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8741 = 9'ha1 == r_count_21_io_out ? io_r_161_b : _GEN_8740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8742 = 9'ha2 == r_count_21_io_out ? io_r_162_b : _GEN_8741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8743 = 9'ha3 == r_count_21_io_out ? io_r_163_b : _GEN_8742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8744 = 9'ha4 == r_count_21_io_out ? io_r_164_b : _GEN_8743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8745 = 9'ha5 == r_count_21_io_out ? io_r_165_b : _GEN_8744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8746 = 9'ha6 == r_count_21_io_out ? io_r_166_b : _GEN_8745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8747 = 9'ha7 == r_count_21_io_out ? io_r_167_b : _GEN_8746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8748 = 9'ha8 == r_count_21_io_out ? io_r_168_b : _GEN_8747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8749 = 9'ha9 == r_count_21_io_out ? io_r_169_b : _GEN_8748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8750 = 9'haa == r_count_21_io_out ? io_r_170_b : _GEN_8749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8751 = 9'hab == r_count_21_io_out ? io_r_171_b : _GEN_8750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8752 = 9'hac == r_count_21_io_out ? io_r_172_b : _GEN_8751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8753 = 9'had == r_count_21_io_out ? io_r_173_b : _GEN_8752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8754 = 9'hae == r_count_21_io_out ? io_r_174_b : _GEN_8753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8755 = 9'haf == r_count_21_io_out ? io_r_175_b : _GEN_8754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8756 = 9'hb0 == r_count_21_io_out ? io_r_176_b : _GEN_8755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8757 = 9'hb1 == r_count_21_io_out ? io_r_177_b : _GEN_8756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8758 = 9'hb2 == r_count_21_io_out ? io_r_178_b : _GEN_8757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8759 = 9'hb3 == r_count_21_io_out ? io_r_179_b : _GEN_8758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8760 = 9'hb4 == r_count_21_io_out ? io_r_180_b : _GEN_8759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8761 = 9'hb5 == r_count_21_io_out ? io_r_181_b : _GEN_8760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8762 = 9'hb6 == r_count_21_io_out ? io_r_182_b : _GEN_8761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8763 = 9'hb7 == r_count_21_io_out ? io_r_183_b : _GEN_8762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8764 = 9'hb8 == r_count_21_io_out ? io_r_184_b : _GEN_8763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8765 = 9'hb9 == r_count_21_io_out ? io_r_185_b : _GEN_8764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8766 = 9'hba == r_count_21_io_out ? io_r_186_b : _GEN_8765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8767 = 9'hbb == r_count_21_io_out ? io_r_187_b : _GEN_8766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8768 = 9'hbc == r_count_21_io_out ? io_r_188_b : _GEN_8767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8769 = 9'hbd == r_count_21_io_out ? io_r_189_b : _GEN_8768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8770 = 9'hbe == r_count_21_io_out ? io_r_190_b : _GEN_8769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8771 = 9'hbf == r_count_21_io_out ? io_r_191_b : _GEN_8770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8772 = 9'hc0 == r_count_21_io_out ? io_r_192_b : _GEN_8771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8773 = 9'hc1 == r_count_21_io_out ? io_r_193_b : _GEN_8772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8774 = 9'hc2 == r_count_21_io_out ? io_r_194_b : _GEN_8773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8775 = 9'hc3 == r_count_21_io_out ? io_r_195_b : _GEN_8774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8776 = 9'hc4 == r_count_21_io_out ? io_r_196_b : _GEN_8775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8777 = 9'hc5 == r_count_21_io_out ? io_r_197_b : _GEN_8776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8778 = 9'hc6 == r_count_21_io_out ? io_r_198_b : _GEN_8777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8779 = 9'hc7 == r_count_21_io_out ? io_r_199_b : _GEN_8778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8780 = 9'hc8 == r_count_21_io_out ? io_r_200_b : _GEN_8779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8781 = 9'hc9 == r_count_21_io_out ? io_r_201_b : _GEN_8780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8782 = 9'hca == r_count_21_io_out ? io_r_202_b : _GEN_8781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8783 = 9'hcb == r_count_21_io_out ? io_r_203_b : _GEN_8782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8784 = 9'hcc == r_count_21_io_out ? io_r_204_b : _GEN_8783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8785 = 9'hcd == r_count_21_io_out ? io_r_205_b : _GEN_8784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8786 = 9'hce == r_count_21_io_out ? io_r_206_b : _GEN_8785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8787 = 9'hcf == r_count_21_io_out ? io_r_207_b : _GEN_8786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8788 = 9'hd0 == r_count_21_io_out ? io_r_208_b : _GEN_8787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8789 = 9'hd1 == r_count_21_io_out ? io_r_209_b : _GEN_8788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8790 = 9'hd2 == r_count_21_io_out ? io_r_210_b : _GEN_8789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8791 = 9'hd3 == r_count_21_io_out ? io_r_211_b : _GEN_8790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8792 = 9'hd4 == r_count_21_io_out ? io_r_212_b : _GEN_8791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8793 = 9'hd5 == r_count_21_io_out ? io_r_213_b : _GEN_8792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8794 = 9'hd6 == r_count_21_io_out ? io_r_214_b : _GEN_8793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8795 = 9'hd7 == r_count_21_io_out ? io_r_215_b : _GEN_8794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8796 = 9'hd8 == r_count_21_io_out ? io_r_216_b : _GEN_8795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8797 = 9'hd9 == r_count_21_io_out ? io_r_217_b : _GEN_8796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8798 = 9'hda == r_count_21_io_out ? io_r_218_b : _GEN_8797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8799 = 9'hdb == r_count_21_io_out ? io_r_219_b : _GEN_8798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8800 = 9'hdc == r_count_21_io_out ? io_r_220_b : _GEN_8799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8801 = 9'hdd == r_count_21_io_out ? io_r_221_b : _GEN_8800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8802 = 9'hde == r_count_21_io_out ? io_r_222_b : _GEN_8801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8803 = 9'hdf == r_count_21_io_out ? io_r_223_b : _GEN_8802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8804 = 9'he0 == r_count_21_io_out ? io_r_224_b : _GEN_8803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8805 = 9'he1 == r_count_21_io_out ? io_r_225_b : _GEN_8804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8806 = 9'he2 == r_count_21_io_out ? io_r_226_b : _GEN_8805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8807 = 9'he3 == r_count_21_io_out ? io_r_227_b : _GEN_8806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8808 = 9'he4 == r_count_21_io_out ? io_r_228_b : _GEN_8807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8809 = 9'he5 == r_count_21_io_out ? io_r_229_b : _GEN_8808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8810 = 9'he6 == r_count_21_io_out ? io_r_230_b : _GEN_8809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8811 = 9'he7 == r_count_21_io_out ? io_r_231_b : _GEN_8810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8812 = 9'he8 == r_count_21_io_out ? io_r_232_b : _GEN_8811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8813 = 9'he9 == r_count_21_io_out ? io_r_233_b : _GEN_8812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8814 = 9'hea == r_count_21_io_out ? io_r_234_b : _GEN_8813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8815 = 9'heb == r_count_21_io_out ? io_r_235_b : _GEN_8814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8816 = 9'hec == r_count_21_io_out ? io_r_236_b : _GEN_8815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8817 = 9'hed == r_count_21_io_out ? io_r_237_b : _GEN_8816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8818 = 9'hee == r_count_21_io_out ? io_r_238_b : _GEN_8817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8819 = 9'hef == r_count_21_io_out ? io_r_239_b : _GEN_8818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8820 = 9'hf0 == r_count_21_io_out ? io_r_240_b : _GEN_8819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8821 = 9'hf1 == r_count_21_io_out ? io_r_241_b : _GEN_8820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8822 = 9'hf2 == r_count_21_io_out ? io_r_242_b : _GEN_8821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8823 = 9'hf3 == r_count_21_io_out ? io_r_243_b : _GEN_8822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8824 = 9'hf4 == r_count_21_io_out ? io_r_244_b : _GEN_8823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8825 = 9'hf5 == r_count_21_io_out ? io_r_245_b : _GEN_8824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8826 = 9'hf6 == r_count_21_io_out ? io_r_246_b : _GEN_8825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8827 = 9'hf7 == r_count_21_io_out ? io_r_247_b : _GEN_8826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8828 = 9'hf8 == r_count_21_io_out ? io_r_248_b : _GEN_8827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8829 = 9'hf9 == r_count_21_io_out ? io_r_249_b : _GEN_8828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8830 = 9'hfa == r_count_21_io_out ? io_r_250_b : _GEN_8829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8831 = 9'hfb == r_count_21_io_out ? io_r_251_b : _GEN_8830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8832 = 9'hfc == r_count_21_io_out ? io_r_252_b : _GEN_8831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8833 = 9'hfd == r_count_21_io_out ? io_r_253_b : _GEN_8832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8834 = 9'hfe == r_count_21_io_out ? io_r_254_b : _GEN_8833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8835 = 9'hff == r_count_21_io_out ? io_r_255_b : _GEN_8834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8836 = 9'h100 == r_count_21_io_out ? io_r_256_b : _GEN_8835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8837 = 9'h101 == r_count_21_io_out ? io_r_257_b : _GEN_8836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8838 = 9'h102 == r_count_21_io_out ? io_r_258_b : _GEN_8837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8839 = 9'h103 == r_count_21_io_out ? io_r_259_b : _GEN_8838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8840 = 9'h104 == r_count_21_io_out ? io_r_260_b : _GEN_8839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8841 = 9'h105 == r_count_21_io_out ? io_r_261_b : _GEN_8840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8842 = 9'h106 == r_count_21_io_out ? io_r_262_b : _GEN_8841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8843 = 9'h107 == r_count_21_io_out ? io_r_263_b : _GEN_8842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8844 = 9'h108 == r_count_21_io_out ? io_r_264_b : _GEN_8843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8845 = 9'h109 == r_count_21_io_out ? io_r_265_b : _GEN_8844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8846 = 9'h10a == r_count_21_io_out ? io_r_266_b : _GEN_8845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8847 = 9'h10b == r_count_21_io_out ? io_r_267_b : _GEN_8846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8848 = 9'h10c == r_count_21_io_out ? io_r_268_b : _GEN_8847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8849 = 9'h10d == r_count_21_io_out ? io_r_269_b : _GEN_8848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8850 = 9'h10e == r_count_21_io_out ? io_r_270_b : _GEN_8849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8851 = 9'h10f == r_count_21_io_out ? io_r_271_b : _GEN_8850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8852 = 9'h110 == r_count_21_io_out ? io_r_272_b : _GEN_8851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8853 = 9'h111 == r_count_21_io_out ? io_r_273_b : _GEN_8852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8854 = 9'h112 == r_count_21_io_out ? io_r_274_b : _GEN_8853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8855 = 9'h113 == r_count_21_io_out ? io_r_275_b : _GEN_8854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8856 = 9'h114 == r_count_21_io_out ? io_r_276_b : _GEN_8855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8857 = 9'h115 == r_count_21_io_out ? io_r_277_b : _GEN_8856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8858 = 9'h116 == r_count_21_io_out ? io_r_278_b : _GEN_8857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8859 = 9'h117 == r_count_21_io_out ? io_r_279_b : _GEN_8858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8860 = 9'h118 == r_count_21_io_out ? io_r_280_b : _GEN_8859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8861 = 9'h119 == r_count_21_io_out ? io_r_281_b : _GEN_8860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8862 = 9'h11a == r_count_21_io_out ? io_r_282_b : _GEN_8861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8863 = 9'h11b == r_count_21_io_out ? io_r_283_b : _GEN_8862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8864 = 9'h11c == r_count_21_io_out ? io_r_284_b : _GEN_8863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8865 = 9'h11d == r_count_21_io_out ? io_r_285_b : _GEN_8864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8866 = 9'h11e == r_count_21_io_out ? io_r_286_b : _GEN_8865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8867 = 9'h11f == r_count_21_io_out ? io_r_287_b : _GEN_8866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8868 = 9'h120 == r_count_21_io_out ? io_r_288_b : _GEN_8867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8869 = 9'h121 == r_count_21_io_out ? io_r_289_b : _GEN_8868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8870 = 9'h122 == r_count_21_io_out ? io_r_290_b : _GEN_8869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8871 = 9'h123 == r_count_21_io_out ? io_r_291_b : _GEN_8870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8872 = 9'h124 == r_count_21_io_out ? io_r_292_b : _GEN_8871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8873 = 9'h125 == r_count_21_io_out ? io_r_293_b : _GEN_8872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8874 = 9'h126 == r_count_21_io_out ? io_r_294_b : _GEN_8873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8875 = 9'h127 == r_count_21_io_out ? io_r_295_b : _GEN_8874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8876 = 9'h128 == r_count_21_io_out ? io_r_296_b : _GEN_8875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8877 = 9'h129 == r_count_21_io_out ? io_r_297_b : _GEN_8876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8878 = 9'h12a == r_count_21_io_out ? io_r_298_b : _GEN_8877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8879 = 9'h12b == r_count_21_io_out ? io_r_299_b : _GEN_8878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8880 = 9'h12c == r_count_21_io_out ? io_r_300_b : _GEN_8879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8881 = 9'h12d == r_count_21_io_out ? io_r_301_b : _GEN_8880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8882 = 9'h12e == r_count_21_io_out ? io_r_302_b : _GEN_8881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8883 = 9'h12f == r_count_21_io_out ? io_r_303_b : _GEN_8882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8884 = 9'h130 == r_count_21_io_out ? io_r_304_b : _GEN_8883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8885 = 9'h131 == r_count_21_io_out ? io_r_305_b : _GEN_8884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8886 = 9'h132 == r_count_21_io_out ? io_r_306_b : _GEN_8885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8887 = 9'h133 == r_count_21_io_out ? io_r_307_b : _GEN_8886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8888 = 9'h134 == r_count_21_io_out ? io_r_308_b : _GEN_8887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8889 = 9'h135 == r_count_21_io_out ? io_r_309_b : _GEN_8888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8890 = 9'h136 == r_count_21_io_out ? io_r_310_b : _GEN_8889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8891 = 9'h137 == r_count_21_io_out ? io_r_311_b : _GEN_8890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8892 = 9'h138 == r_count_21_io_out ? io_r_312_b : _GEN_8891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8893 = 9'h139 == r_count_21_io_out ? io_r_313_b : _GEN_8892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8894 = 9'h13a == r_count_21_io_out ? io_r_314_b : _GEN_8893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8895 = 9'h13b == r_count_21_io_out ? io_r_315_b : _GEN_8894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8896 = 9'h13c == r_count_21_io_out ? io_r_316_b : _GEN_8895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8897 = 9'h13d == r_count_21_io_out ? io_r_317_b : _GEN_8896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8898 = 9'h13e == r_count_21_io_out ? io_r_318_b : _GEN_8897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8899 = 9'h13f == r_count_21_io_out ? io_r_319_b : _GEN_8898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8900 = 9'h140 == r_count_21_io_out ? io_r_320_b : _GEN_8899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8901 = 9'h141 == r_count_21_io_out ? io_r_321_b : _GEN_8900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8902 = 9'h142 == r_count_21_io_out ? io_r_322_b : _GEN_8901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8903 = 9'h143 == r_count_21_io_out ? io_r_323_b : _GEN_8902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8904 = 9'h144 == r_count_21_io_out ? io_r_324_b : _GEN_8903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8905 = 9'h145 == r_count_21_io_out ? io_r_325_b : _GEN_8904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8906 = 9'h146 == r_count_21_io_out ? io_r_326_b : _GEN_8905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8907 = 9'h147 == r_count_21_io_out ? io_r_327_b : _GEN_8906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8908 = 9'h148 == r_count_21_io_out ? io_r_328_b : _GEN_8907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8909 = 9'h149 == r_count_21_io_out ? io_r_329_b : _GEN_8908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8910 = 9'h14a == r_count_21_io_out ? io_r_330_b : _GEN_8909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8911 = 9'h14b == r_count_21_io_out ? io_r_331_b : _GEN_8910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8912 = 9'h14c == r_count_21_io_out ? io_r_332_b : _GEN_8911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8913 = 9'h14d == r_count_21_io_out ? io_r_333_b : _GEN_8912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8914 = 9'h14e == r_count_21_io_out ? io_r_334_b : _GEN_8913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8915 = 9'h14f == r_count_21_io_out ? io_r_335_b : _GEN_8914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8916 = 9'h150 == r_count_21_io_out ? io_r_336_b : _GEN_8915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8917 = 9'h151 == r_count_21_io_out ? io_r_337_b : _GEN_8916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8918 = 9'h152 == r_count_21_io_out ? io_r_338_b : _GEN_8917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8919 = 9'h153 == r_count_21_io_out ? io_r_339_b : _GEN_8918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8920 = 9'h154 == r_count_21_io_out ? io_r_340_b : _GEN_8919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8921 = 9'h155 == r_count_21_io_out ? io_r_341_b : _GEN_8920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8922 = 9'h156 == r_count_21_io_out ? io_r_342_b : _GEN_8921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8923 = 9'h157 == r_count_21_io_out ? io_r_343_b : _GEN_8922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8924 = 9'h158 == r_count_21_io_out ? io_r_344_b : _GEN_8923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8925 = 9'h159 == r_count_21_io_out ? io_r_345_b : _GEN_8924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8926 = 9'h15a == r_count_21_io_out ? io_r_346_b : _GEN_8925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8927 = 9'h15b == r_count_21_io_out ? io_r_347_b : _GEN_8926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8928 = 9'h15c == r_count_21_io_out ? io_r_348_b : _GEN_8927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8929 = 9'h15d == r_count_21_io_out ? io_r_349_b : _GEN_8928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8930 = 9'h15e == r_count_21_io_out ? io_r_350_b : _GEN_8929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8931 = 9'h15f == r_count_21_io_out ? io_r_351_b : _GEN_8930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8932 = 9'h160 == r_count_21_io_out ? io_r_352_b : _GEN_8931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8933 = 9'h161 == r_count_21_io_out ? io_r_353_b : _GEN_8932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8934 = 9'h162 == r_count_21_io_out ? io_r_354_b : _GEN_8933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8935 = 9'h163 == r_count_21_io_out ? io_r_355_b : _GEN_8934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8936 = 9'h164 == r_count_21_io_out ? io_r_356_b : _GEN_8935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8937 = 9'h165 == r_count_21_io_out ? io_r_357_b : _GEN_8936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8938 = 9'h166 == r_count_21_io_out ? io_r_358_b : _GEN_8937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8939 = 9'h167 == r_count_21_io_out ? io_r_359_b : _GEN_8938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8940 = 9'h168 == r_count_21_io_out ? io_r_360_b : _GEN_8939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8941 = 9'h169 == r_count_21_io_out ? io_r_361_b : _GEN_8940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8942 = 9'h16a == r_count_21_io_out ? io_r_362_b : _GEN_8941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8943 = 9'h16b == r_count_21_io_out ? io_r_363_b : _GEN_8942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8944 = 9'h16c == r_count_21_io_out ? io_r_364_b : _GEN_8943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8945 = 9'h16d == r_count_21_io_out ? io_r_365_b : _GEN_8944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8946 = 9'h16e == r_count_21_io_out ? io_r_366_b : _GEN_8945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8947 = 9'h16f == r_count_21_io_out ? io_r_367_b : _GEN_8946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8948 = 9'h170 == r_count_21_io_out ? io_r_368_b : _GEN_8947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8949 = 9'h171 == r_count_21_io_out ? io_r_369_b : _GEN_8948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8950 = 9'h172 == r_count_21_io_out ? io_r_370_b : _GEN_8949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8951 = 9'h173 == r_count_21_io_out ? io_r_371_b : _GEN_8950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8952 = 9'h174 == r_count_21_io_out ? io_r_372_b : _GEN_8951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8953 = 9'h175 == r_count_21_io_out ? io_r_373_b : _GEN_8952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8954 = 9'h176 == r_count_21_io_out ? io_r_374_b : _GEN_8953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8955 = 9'h177 == r_count_21_io_out ? io_r_375_b : _GEN_8954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8956 = 9'h178 == r_count_21_io_out ? io_r_376_b : _GEN_8955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8957 = 9'h179 == r_count_21_io_out ? io_r_377_b : _GEN_8956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8958 = 9'h17a == r_count_21_io_out ? io_r_378_b : _GEN_8957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8959 = 9'h17b == r_count_21_io_out ? io_r_379_b : _GEN_8958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8960 = 9'h17c == r_count_21_io_out ? io_r_380_b : _GEN_8959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8961 = 9'h17d == r_count_21_io_out ? io_r_381_b : _GEN_8960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8962 = 9'h17e == r_count_21_io_out ? io_r_382_b : _GEN_8961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8963 = 9'h17f == r_count_21_io_out ? io_r_383_b : _GEN_8962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8964 = 9'h180 == r_count_21_io_out ? io_r_384_b : _GEN_8963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8965 = 9'h181 == r_count_21_io_out ? io_r_385_b : _GEN_8964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8966 = 9'h182 == r_count_21_io_out ? io_r_386_b : _GEN_8965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8967 = 9'h183 == r_count_21_io_out ? io_r_387_b : _GEN_8966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8968 = 9'h184 == r_count_21_io_out ? io_r_388_b : _GEN_8967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8969 = 9'h185 == r_count_21_io_out ? io_r_389_b : _GEN_8968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8970 = 9'h186 == r_count_21_io_out ? io_r_390_b : _GEN_8969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8971 = 9'h187 == r_count_21_io_out ? io_r_391_b : _GEN_8970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8972 = 9'h188 == r_count_21_io_out ? io_r_392_b : _GEN_8971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8973 = 9'h189 == r_count_21_io_out ? io_r_393_b : _GEN_8972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8974 = 9'h18a == r_count_21_io_out ? io_r_394_b : _GEN_8973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8975 = 9'h18b == r_count_21_io_out ? io_r_395_b : _GEN_8974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8976 = 9'h18c == r_count_21_io_out ? io_r_396_b : _GEN_8975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8977 = 9'h18d == r_count_21_io_out ? io_r_397_b : _GEN_8976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8978 = 9'h18e == r_count_21_io_out ? io_r_398_b : _GEN_8977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8981 = 9'h1 == r_count_22_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8982 = 9'h2 == r_count_22_io_out ? io_r_2_b : _GEN_8981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8983 = 9'h3 == r_count_22_io_out ? io_r_3_b : _GEN_8982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8984 = 9'h4 == r_count_22_io_out ? io_r_4_b : _GEN_8983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8985 = 9'h5 == r_count_22_io_out ? io_r_5_b : _GEN_8984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8986 = 9'h6 == r_count_22_io_out ? io_r_6_b : _GEN_8985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8987 = 9'h7 == r_count_22_io_out ? io_r_7_b : _GEN_8986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8988 = 9'h8 == r_count_22_io_out ? io_r_8_b : _GEN_8987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8989 = 9'h9 == r_count_22_io_out ? io_r_9_b : _GEN_8988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8990 = 9'ha == r_count_22_io_out ? io_r_10_b : _GEN_8989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8991 = 9'hb == r_count_22_io_out ? io_r_11_b : _GEN_8990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8992 = 9'hc == r_count_22_io_out ? io_r_12_b : _GEN_8991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8993 = 9'hd == r_count_22_io_out ? io_r_13_b : _GEN_8992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8994 = 9'he == r_count_22_io_out ? io_r_14_b : _GEN_8993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8995 = 9'hf == r_count_22_io_out ? io_r_15_b : _GEN_8994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8996 = 9'h10 == r_count_22_io_out ? io_r_16_b : _GEN_8995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8997 = 9'h11 == r_count_22_io_out ? io_r_17_b : _GEN_8996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8998 = 9'h12 == r_count_22_io_out ? io_r_18_b : _GEN_8997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8999 = 9'h13 == r_count_22_io_out ? io_r_19_b : _GEN_8998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9000 = 9'h14 == r_count_22_io_out ? io_r_20_b : _GEN_8999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9001 = 9'h15 == r_count_22_io_out ? io_r_21_b : _GEN_9000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9002 = 9'h16 == r_count_22_io_out ? io_r_22_b : _GEN_9001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9003 = 9'h17 == r_count_22_io_out ? io_r_23_b : _GEN_9002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9004 = 9'h18 == r_count_22_io_out ? io_r_24_b : _GEN_9003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9005 = 9'h19 == r_count_22_io_out ? io_r_25_b : _GEN_9004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9006 = 9'h1a == r_count_22_io_out ? io_r_26_b : _GEN_9005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9007 = 9'h1b == r_count_22_io_out ? io_r_27_b : _GEN_9006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9008 = 9'h1c == r_count_22_io_out ? io_r_28_b : _GEN_9007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9009 = 9'h1d == r_count_22_io_out ? io_r_29_b : _GEN_9008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9010 = 9'h1e == r_count_22_io_out ? io_r_30_b : _GEN_9009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9011 = 9'h1f == r_count_22_io_out ? io_r_31_b : _GEN_9010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9012 = 9'h20 == r_count_22_io_out ? io_r_32_b : _GEN_9011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9013 = 9'h21 == r_count_22_io_out ? io_r_33_b : _GEN_9012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9014 = 9'h22 == r_count_22_io_out ? io_r_34_b : _GEN_9013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9015 = 9'h23 == r_count_22_io_out ? io_r_35_b : _GEN_9014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9016 = 9'h24 == r_count_22_io_out ? io_r_36_b : _GEN_9015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9017 = 9'h25 == r_count_22_io_out ? io_r_37_b : _GEN_9016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9018 = 9'h26 == r_count_22_io_out ? io_r_38_b : _GEN_9017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9019 = 9'h27 == r_count_22_io_out ? io_r_39_b : _GEN_9018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9020 = 9'h28 == r_count_22_io_out ? io_r_40_b : _GEN_9019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9021 = 9'h29 == r_count_22_io_out ? io_r_41_b : _GEN_9020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9022 = 9'h2a == r_count_22_io_out ? io_r_42_b : _GEN_9021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9023 = 9'h2b == r_count_22_io_out ? io_r_43_b : _GEN_9022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9024 = 9'h2c == r_count_22_io_out ? io_r_44_b : _GEN_9023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9025 = 9'h2d == r_count_22_io_out ? io_r_45_b : _GEN_9024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9026 = 9'h2e == r_count_22_io_out ? io_r_46_b : _GEN_9025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9027 = 9'h2f == r_count_22_io_out ? io_r_47_b : _GEN_9026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9028 = 9'h30 == r_count_22_io_out ? io_r_48_b : _GEN_9027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9029 = 9'h31 == r_count_22_io_out ? io_r_49_b : _GEN_9028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9030 = 9'h32 == r_count_22_io_out ? io_r_50_b : _GEN_9029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9031 = 9'h33 == r_count_22_io_out ? io_r_51_b : _GEN_9030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9032 = 9'h34 == r_count_22_io_out ? io_r_52_b : _GEN_9031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9033 = 9'h35 == r_count_22_io_out ? io_r_53_b : _GEN_9032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9034 = 9'h36 == r_count_22_io_out ? io_r_54_b : _GEN_9033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9035 = 9'h37 == r_count_22_io_out ? io_r_55_b : _GEN_9034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9036 = 9'h38 == r_count_22_io_out ? io_r_56_b : _GEN_9035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9037 = 9'h39 == r_count_22_io_out ? io_r_57_b : _GEN_9036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9038 = 9'h3a == r_count_22_io_out ? io_r_58_b : _GEN_9037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9039 = 9'h3b == r_count_22_io_out ? io_r_59_b : _GEN_9038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9040 = 9'h3c == r_count_22_io_out ? io_r_60_b : _GEN_9039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9041 = 9'h3d == r_count_22_io_out ? io_r_61_b : _GEN_9040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9042 = 9'h3e == r_count_22_io_out ? io_r_62_b : _GEN_9041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9043 = 9'h3f == r_count_22_io_out ? io_r_63_b : _GEN_9042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9044 = 9'h40 == r_count_22_io_out ? io_r_64_b : _GEN_9043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9045 = 9'h41 == r_count_22_io_out ? io_r_65_b : _GEN_9044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9046 = 9'h42 == r_count_22_io_out ? io_r_66_b : _GEN_9045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9047 = 9'h43 == r_count_22_io_out ? io_r_67_b : _GEN_9046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9048 = 9'h44 == r_count_22_io_out ? io_r_68_b : _GEN_9047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9049 = 9'h45 == r_count_22_io_out ? io_r_69_b : _GEN_9048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9050 = 9'h46 == r_count_22_io_out ? io_r_70_b : _GEN_9049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9051 = 9'h47 == r_count_22_io_out ? io_r_71_b : _GEN_9050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9052 = 9'h48 == r_count_22_io_out ? io_r_72_b : _GEN_9051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9053 = 9'h49 == r_count_22_io_out ? io_r_73_b : _GEN_9052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9054 = 9'h4a == r_count_22_io_out ? io_r_74_b : _GEN_9053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9055 = 9'h4b == r_count_22_io_out ? io_r_75_b : _GEN_9054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9056 = 9'h4c == r_count_22_io_out ? io_r_76_b : _GEN_9055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9057 = 9'h4d == r_count_22_io_out ? io_r_77_b : _GEN_9056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9058 = 9'h4e == r_count_22_io_out ? io_r_78_b : _GEN_9057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9059 = 9'h4f == r_count_22_io_out ? io_r_79_b : _GEN_9058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9060 = 9'h50 == r_count_22_io_out ? io_r_80_b : _GEN_9059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9061 = 9'h51 == r_count_22_io_out ? io_r_81_b : _GEN_9060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9062 = 9'h52 == r_count_22_io_out ? io_r_82_b : _GEN_9061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9063 = 9'h53 == r_count_22_io_out ? io_r_83_b : _GEN_9062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9064 = 9'h54 == r_count_22_io_out ? io_r_84_b : _GEN_9063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9065 = 9'h55 == r_count_22_io_out ? io_r_85_b : _GEN_9064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9066 = 9'h56 == r_count_22_io_out ? io_r_86_b : _GEN_9065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9067 = 9'h57 == r_count_22_io_out ? io_r_87_b : _GEN_9066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9068 = 9'h58 == r_count_22_io_out ? io_r_88_b : _GEN_9067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9069 = 9'h59 == r_count_22_io_out ? io_r_89_b : _GEN_9068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9070 = 9'h5a == r_count_22_io_out ? io_r_90_b : _GEN_9069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9071 = 9'h5b == r_count_22_io_out ? io_r_91_b : _GEN_9070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9072 = 9'h5c == r_count_22_io_out ? io_r_92_b : _GEN_9071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9073 = 9'h5d == r_count_22_io_out ? io_r_93_b : _GEN_9072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9074 = 9'h5e == r_count_22_io_out ? io_r_94_b : _GEN_9073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9075 = 9'h5f == r_count_22_io_out ? io_r_95_b : _GEN_9074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9076 = 9'h60 == r_count_22_io_out ? io_r_96_b : _GEN_9075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9077 = 9'h61 == r_count_22_io_out ? io_r_97_b : _GEN_9076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9078 = 9'h62 == r_count_22_io_out ? io_r_98_b : _GEN_9077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9079 = 9'h63 == r_count_22_io_out ? io_r_99_b : _GEN_9078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9080 = 9'h64 == r_count_22_io_out ? io_r_100_b : _GEN_9079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9081 = 9'h65 == r_count_22_io_out ? io_r_101_b : _GEN_9080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9082 = 9'h66 == r_count_22_io_out ? io_r_102_b : _GEN_9081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9083 = 9'h67 == r_count_22_io_out ? io_r_103_b : _GEN_9082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9084 = 9'h68 == r_count_22_io_out ? io_r_104_b : _GEN_9083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9085 = 9'h69 == r_count_22_io_out ? io_r_105_b : _GEN_9084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9086 = 9'h6a == r_count_22_io_out ? io_r_106_b : _GEN_9085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9087 = 9'h6b == r_count_22_io_out ? io_r_107_b : _GEN_9086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9088 = 9'h6c == r_count_22_io_out ? io_r_108_b : _GEN_9087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9089 = 9'h6d == r_count_22_io_out ? io_r_109_b : _GEN_9088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9090 = 9'h6e == r_count_22_io_out ? io_r_110_b : _GEN_9089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9091 = 9'h6f == r_count_22_io_out ? io_r_111_b : _GEN_9090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9092 = 9'h70 == r_count_22_io_out ? io_r_112_b : _GEN_9091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9093 = 9'h71 == r_count_22_io_out ? io_r_113_b : _GEN_9092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9094 = 9'h72 == r_count_22_io_out ? io_r_114_b : _GEN_9093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9095 = 9'h73 == r_count_22_io_out ? io_r_115_b : _GEN_9094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9096 = 9'h74 == r_count_22_io_out ? io_r_116_b : _GEN_9095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9097 = 9'h75 == r_count_22_io_out ? io_r_117_b : _GEN_9096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9098 = 9'h76 == r_count_22_io_out ? io_r_118_b : _GEN_9097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9099 = 9'h77 == r_count_22_io_out ? io_r_119_b : _GEN_9098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9100 = 9'h78 == r_count_22_io_out ? io_r_120_b : _GEN_9099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9101 = 9'h79 == r_count_22_io_out ? io_r_121_b : _GEN_9100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9102 = 9'h7a == r_count_22_io_out ? io_r_122_b : _GEN_9101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9103 = 9'h7b == r_count_22_io_out ? io_r_123_b : _GEN_9102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9104 = 9'h7c == r_count_22_io_out ? io_r_124_b : _GEN_9103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9105 = 9'h7d == r_count_22_io_out ? io_r_125_b : _GEN_9104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9106 = 9'h7e == r_count_22_io_out ? io_r_126_b : _GEN_9105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9107 = 9'h7f == r_count_22_io_out ? io_r_127_b : _GEN_9106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9108 = 9'h80 == r_count_22_io_out ? io_r_128_b : _GEN_9107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9109 = 9'h81 == r_count_22_io_out ? io_r_129_b : _GEN_9108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9110 = 9'h82 == r_count_22_io_out ? io_r_130_b : _GEN_9109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9111 = 9'h83 == r_count_22_io_out ? io_r_131_b : _GEN_9110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9112 = 9'h84 == r_count_22_io_out ? io_r_132_b : _GEN_9111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9113 = 9'h85 == r_count_22_io_out ? io_r_133_b : _GEN_9112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9114 = 9'h86 == r_count_22_io_out ? io_r_134_b : _GEN_9113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9115 = 9'h87 == r_count_22_io_out ? io_r_135_b : _GEN_9114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9116 = 9'h88 == r_count_22_io_out ? io_r_136_b : _GEN_9115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9117 = 9'h89 == r_count_22_io_out ? io_r_137_b : _GEN_9116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9118 = 9'h8a == r_count_22_io_out ? io_r_138_b : _GEN_9117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9119 = 9'h8b == r_count_22_io_out ? io_r_139_b : _GEN_9118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9120 = 9'h8c == r_count_22_io_out ? io_r_140_b : _GEN_9119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9121 = 9'h8d == r_count_22_io_out ? io_r_141_b : _GEN_9120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9122 = 9'h8e == r_count_22_io_out ? io_r_142_b : _GEN_9121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9123 = 9'h8f == r_count_22_io_out ? io_r_143_b : _GEN_9122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9124 = 9'h90 == r_count_22_io_out ? io_r_144_b : _GEN_9123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9125 = 9'h91 == r_count_22_io_out ? io_r_145_b : _GEN_9124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9126 = 9'h92 == r_count_22_io_out ? io_r_146_b : _GEN_9125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9127 = 9'h93 == r_count_22_io_out ? io_r_147_b : _GEN_9126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9128 = 9'h94 == r_count_22_io_out ? io_r_148_b : _GEN_9127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9129 = 9'h95 == r_count_22_io_out ? io_r_149_b : _GEN_9128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9130 = 9'h96 == r_count_22_io_out ? io_r_150_b : _GEN_9129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9131 = 9'h97 == r_count_22_io_out ? io_r_151_b : _GEN_9130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9132 = 9'h98 == r_count_22_io_out ? io_r_152_b : _GEN_9131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9133 = 9'h99 == r_count_22_io_out ? io_r_153_b : _GEN_9132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9134 = 9'h9a == r_count_22_io_out ? io_r_154_b : _GEN_9133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9135 = 9'h9b == r_count_22_io_out ? io_r_155_b : _GEN_9134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9136 = 9'h9c == r_count_22_io_out ? io_r_156_b : _GEN_9135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9137 = 9'h9d == r_count_22_io_out ? io_r_157_b : _GEN_9136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9138 = 9'h9e == r_count_22_io_out ? io_r_158_b : _GEN_9137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9139 = 9'h9f == r_count_22_io_out ? io_r_159_b : _GEN_9138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9140 = 9'ha0 == r_count_22_io_out ? io_r_160_b : _GEN_9139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9141 = 9'ha1 == r_count_22_io_out ? io_r_161_b : _GEN_9140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9142 = 9'ha2 == r_count_22_io_out ? io_r_162_b : _GEN_9141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9143 = 9'ha3 == r_count_22_io_out ? io_r_163_b : _GEN_9142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9144 = 9'ha4 == r_count_22_io_out ? io_r_164_b : _GEN_9143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9145 = 9'ha5 == r_count_22_io_out ? io_r_165_b : _GEN_9144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9146 = 9'ha6 == r_count_22_io_out ? io_r_166_b : _GEN_9145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9147 = 9'ha7 == r_count_22_io_out ? io_r_167_b : _GEN_9146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9148 = 9'ha8 == r_count_22_io_out ? io_r_168_b : _GEN_9147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9149 = 9'ha9 == r_count_22_io_out ? io_r_169_b : _GEN_9148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9150 = 9'haa == r_count_22_io_out ? io_r_170_b : _GEN_9149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9151 = 9'hab == r_count_22_io_out ? io_r_171_b : _GEN_9150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9152 = 9'hac == r_count_22_io_out ? io_r_172_b : _GEN_9151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9153 = 9'had == r_count_22_io_out ? io_r_173_b : _GEN_9152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9154 = 9'hae == r_count_22_io_out ? io_r_174_b : _GEN_9153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9155 = 9'haf == r_count_22_io_out ? io_r_175_b : _GEN_9154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9156 = 9'hb0 == r_count_22_io_out ? io_r_176_b : _GEN_9155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9157 = 9'hb1 == r_count_22_io_out ? io_r_177_b : _GEN_9156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9158 = 9'hb2 == r_count_22_io_out ? io_r_178_b : _GEN_9157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9159 = 9'hb3 == r_count_22_io_out ? io_r_179_b : _GEN_9158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9160 = 9'hb4 == r_count_22_io_out ? io_r_180_b : _GEN_9159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9161 = 9'hb5 == r_count_22_io_out ? io_r_181_b : _GEN_9160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9162 = 9'hb6 == r_count_22_io_out ? io_r_182_b : _GEN_9161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9163 = 9'hb7 == r_count_22_io_out ? io_r_183_b : _GEN_9162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9164 = 9'hb8 == r_count_22_io_out ? io_r_184_b : _GEN_9163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9165 = 9'hb9 == r_count_22_io_out ? io_r_185_b : _GEN_9164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9166 = 9'hba == r_count_22_io_out ? io_r_186_b : _GEN_9165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9167 = 9'hbb == r_count_22_io_out ? io_r_187_b : _GEN_9166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9168 = 9'hbc == r_count_22_io_out ? io_r_188_b : _GEN_9167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9169 = 9'hbd == r_count_22_io_out ? io_r_189_b : _GEN_9168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9170 = 9'hbe == r_count_22_io_out ? io_r_190_b : _GEN_9169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9171 = 9'hbf == r_count_22_io_out ? io_r_191_b : _GEN_9170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9172 = 9'hc0 == r_count_22_io_out ? io_r_192_b : _GEN_9171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9173 = 9'hc1 == r_count_22_io_out ? io_r_193_b : _GEN_9172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9174 = 9'hc2 == r_count_22_io_out ? io_r_194_b : _GEN_9173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9175 = 9'hc3 == r_count_22_io_out ? io_r_195_b : _GEN_9174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9176 = 9'hc4 == r_count_22_io_out ? io_r_196_b : _GEN_9175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9177 = 9'hc5 == r_count_22_io_out ? io_r_197_b : _GEN_9176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9178 = 9'hc6 == r_count_22_io_out ? io_r_198_b : _GEN_9177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9179 = 9'hc7 == r_count_22_io_out ? io_r_199_b : _GEN_9178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9180 = 9'hc8 == r_count_22_io_out ? io_r_200_b : _GEN_9179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9181 = 9'hc9 == r_count_22_io_out ? io_r_201_b : _GEN_9180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9182 = 9'hca == r_count_22_io_out ? io_r_202_b : _GEN_9181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9183 = 9'hcb == r_count_22_io_out ? io_r_203_b : _GEN_9182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9184 = 9'hcc == r_count_22_io_out ? io_r_204_b : _GEN_9183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9185 = 9'hcd == r_count_22_io_out ? io_r_205_b : _GEN_9184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9186 = 9'hce == r_count_22_io_out ? io_r_206_b : _GEN_9185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9187 = 9'hcf == r_count_22_io_out ? io_r_207_b : _GEN_9186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9188 = 9'hd0 == r_count_22_io_out ? io_r_208_b : _GEN_9187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9189 = 9'hd1 == r_count_22_io_out ? io_r_209_b : _GEN_9188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9190 = 9'hd2 == r_count_22_io_out ? io_r_210_b : _GEN_9189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9191 = 9'hd3 == r_count_22_io_out ? io_r_211_b : _GEN_9190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9192 = 9'hd4 == r_count_22_io_out ? io_r_212_b : _GEN_9191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9193 = 9'hd5 == r_count_22_io_out ? io_r_213_b : _GEN_9192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9194 = 9'hd6 == r_count_22_io_out ? io_r_214_b : _GEN_9193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9195 = 9'hd7 == r_count_22_io_out ? io_r_215_b : _GEN_9194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9196 = 9'hd8 == r_count_22_io_out ? io_r_216_b : _GEN_9195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9197 = 9'hd9 == r_count_22_io_out ? io_r_217_b : _GEN_9196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9198 = 9'hda == r_count_22_io_out ? io_r_218_b : _GEN_9197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9199 = 9'hdb == r_count_22_io_out ? io_r_219_b : _GEN_9198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9200 = 9'hdc == r_count_22_io_out ? io_r_220_b : _GEN_9199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9201 = 9'hdd == r_count_22_io_out ? io_r_221_b : _GEN_9200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9202 = 9'hde == r_count_22_io_out ? io_r_222_b : _GEN_9201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9203 = 9'hdf == r_count_22_io_out ? io_r_223_b : _GEN_9202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9204 = 9'he0 == r_count_22_io_out ? io_r_224_b : _GEN_9203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9205 = 9'he1 == r_count_22_io_out ? io_r_225_b : _GEN_9204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9206 = 9'he2 == r_count_22_io_out ? io_r_226_b : _GEN_9205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9207 = 9'he3 == r_count_22_io_out ? io_r_227_b : _GEN_9206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9208 = 9'he4 == r_count_22_io_out ? io_r_228_b : _GEN_9207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9209 = 9'he5 == r_count_22_io_out ? io_r_229_b : _GEN_9208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9210 = 9'he6 == r_count_22_io_out ? io_r_230_b : _GEN_9209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9211 = 9'he7 == r_count_22_io_out ? io_r_231_b : _GEN_9210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9212 = 9'he8 == r_count_22_io_out ? io_r_232_b : _GEN_9211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9213 = 9'he9 == r_count_22_io_out ? io_r_233_b : _GEN_9212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9214 = 9'hea == r_count_22_io_out ? io_r_234_b : _GEN_9213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9215 = 9'heb == r_count_22_io_out ? io_r_235_b : _GEN_9214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9216 = 9'hec == r_count_22_io_out ? io_r_236_b : _GEN_9215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9217 = 9'hed == r_count_22_io_out ? io_r_237_b : _GEN_9216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9218 = 9'hee == r_count_22_io_out ? io_r_238_b : _GEN_9217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9219 = 9'hef == r_count_22_io_out ? io_r_239_b : _GEN_9218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9220 = 9'hf0 == r_count_22_io_out ? io_r_240_b : _GEN_9219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9221 = 9'hf1 == r_count_22_io_out ? io_r_241_b : _GEN_9220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9222 = 9'hf2 == r_count_22_io_out ? io_r_242_b : _GEN_9221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9223 = 9'hf3 == r_count_22_io_out ? io_r_243_b : _GEN_9222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9224 = 9'hf4 == r_count_22_io_out ? io_r_244_b : _GEN_9223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9225 = 9'hf5 == r_count_22_io_out ? io_r_245_b : _GEN_9224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9226 = 9'hf6 == r_count_22_io_out ? io_r_246_b : _GEN_9225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9227 = 9'hf7 == r_count_22_io_out ? io_r_247_b : _GEN_9226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9228 = 9'hf8 == r_count_22_io_out ? io_r_248_b : _GEN_9227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9229 = 9'hf9 == r_count_22_io_out ? io_r_249_b : _GEN_9228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9230 = 9'hfa == r_count_22_io_out ? io_r_250_b : _GEN_9229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9231 = 9'hfb == r_count_22_io_out ? io_r_251_b : _GEN_9230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9232 = 9'hfc == r_count_22_io_out ? io_r_252_b : _GEN_9231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9233 = 9'hfd == r_count_22_io_out ? io_r_253_b : _GEN_9232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9234 = 9'hfe == r_count_22_io_out ? io_r_254_b : _GEN_9233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9235 = 9'hff == r_count_22_io_out ? io_r_255_b : _GEN_9234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9236 = 9'h100 == r_count_22_io_out ? io_r_256_b : _GEN_9235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9237 = 9'h101 == r_count_22_io_out ? io_r_257_b : _GEN_9236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9238 = 9'h102 == r_count_22_io_out ? io_r_258_b : _GEN_9237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9239 = 9'h103 == r_count_22_io_out ? io_r_259_b : _GEN_9238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9240 = 9'h104 == r_count_22_io_out ? io_r_260_b : _GEN_9239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9241 = 9'h105 == r_count_22_io_out ? io_r_261_b : _GEN_9240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9242 = 9'h106 == r_count_22_io_out ? io_r_262_b : _GEN_9241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9243 = 9'h107 == r_count_22_io_out ? io_r_263_b : _GEN_9242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9244 = 9'h108 == r_count_22_io_out ? io_r_264_b : _GEN_9243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9245 = 9'h109 == r_count_22_io_out ? io_r_265_b : _GEN_9244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9246 = 9'h10a == r_count_22_io_out ? io_r_266_b : _GEN_9245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9247 = 9'h10b == r_count_22_io_out ? io_r_267_b : _GEN_9246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9248 = 9'h10c == r_count_22_io_out ? io_r_268_b : _GEN_9247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9249 = 9'h10d == r_count_22_io_out ? io_r_269_b : _GEN_9248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9250 = 9'h10e == r_count_22_io_out ? io_r_270_b : _GEN_9249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9251 = 9'h10f == r_count_22_io_out ? io_r_271_b : _GEN_9250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9252 = 9'h110 == r_count_22_io_out ? io_r_272_b : _GEN_9251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9253 = 9'h111 == r_count_22_io_out ? io_r_273_b : _GEN_9252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9254 = 9'h112 == r_count_22_io_out ? io_r_274_b : _GEN_9253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9255 = 9'h113 == r_count_22_io_out ? io_r_275_b : _GEN_9254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9256 = 9'h114 == r_count_22_io_out ? io_r_276_b : _GEN_9255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9257 = 9'h115 == r_count_22_io_out ? io_r_277_b : _GEN_9256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9258 = 9'h116 == r_count_22_io_out ? io_r_278_b : _GEN_9257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9259 = 9'h117 == r_count_22_io_out ? io_r_279_b : _GEN_9258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9260 = 9'h118 == r_count_22_io_out ? io_r_280_b : _GEN_9259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9261 = 9'h119 == r_count_22_io_out ? io_r_281_b : _GEN_9260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9262 = 9'h11a == r_count_22_io_out ? io_r_282_b : _GEN_9261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9263 = 9'h11b == r_count_22_io_out ? io_r_283_b : _GEN_9262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9264 = 9'h11c == r_count_22_io_out ? io_r_284_b : _GEN_9263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9265 = 9'h11d == r_count_22_io_out ? io_r_285_b : _GEN_9264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9266 = 9'h11e == r_count_22_io_out ? io_r_286_b : _GEN_9265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9267 = 9'h11f == r_count_22_io_out ? io_r_287_b : _GEN_9266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9268 = 9'h120 == r_count_22_io_out ? io_r_288_b : _GEN_9267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9269 = 9'h121 == r_count_22_io_out ? io_r_289_b : _GEN_9268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9270 = 9'h122 == r_count_22_io_out ? io_r_290_b : _GEN_9269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9271 = 9'h123 == r_count_22_io_out ? io_r_291_b : _GEN_9270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9272 = 9'h124 == r_count_22_io_out ? io_r_292_b : _GEN_9271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9273 = 9'h125 == r_count_22_io_out ? io_r_293_b : _GEN_9272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9274 = 9'h126 == r_count_22_io_out ? io_r_294_b : _GEN_9273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9275 = 9'h127 == r_count_22_io_out ? io_r_295_b : _GEN_9274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9276 = 9'h128 == r_count_22_io_out ? io_r_296_b : _GEN_9275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9277 = 9'h129 == r_count_22_io_out ? io_r_297_b : _GEN_9276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9278 = 9'h12a == r_count_22_io_out ? io_r_298_b : _GEN_9277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9279 = 9'h12b == r_count_22_io_out ? io_r_299_b : _GEN_9278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9280 = 9'h12c == r_count_22_io_out ? io_r_300_b : _GEN_9279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9281 = 9'h12d == r_count_22_io_out ? io_r_301_b : _GEN_9280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9282 = 9'h12e == r_count_22_io_out ? io_r_302_b : _GEN_9281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9283 = 9'h12f == r_count_22_io_out ? io_r_303_b : _GEN_9282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9284 = 9'h130 == r_count_22_io_out ? io_r_304_b : _GEN_9283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9285 = 9'h131 == r_count_22_io_out ? io_r_305_b : _GEN_9284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9286 = 9'h132 == r_count_22_io_out ? io_r_306_b : _GEN_9285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9287 = 9'h133 == r_count_22_io_out ? io_r_307_b : _GEN_9286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9288 = 9'h134 == r_count_22_io_out ? io_r_308_b : _GEN_9287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9289 = 9'h135 == r_count_22_io_out ? io_r_309_b : _GEN_9288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9290 = 9'h136 == r_count_22_io_out ? io_r_310_b : _GEN_9289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9291 = 9'h137 == r_count_22_io_out ? io_r_311_b : _GEN_9290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9292 = 9'h138 == r_count_22_io_out ? io_r_312_b : _GEN_9291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9293 = 9'h139 == r_count_22_io_out ? io_r_313_b : _GEN_9292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9294 = 9'h13a == r_count_22_io_out ? io_r_314_b : _GEN_9293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9295 = 9'h13b == r_count_22_io_out ? io_r_315_b : _GEN_9294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9296 = 9'h13c == r_count_22_io_out ? io_r_316_b : _GEN_9295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9297 = 9'h13d == r_count_22_io_out ? io_r_317_b : _GEN_9296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9298 = 9'h13e == r_count_22_io_out ? io_r_318_b : _GEN_9297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9299 = 9'h13f == r_count_22_io_out ? io_r_319_b : _GEN_9298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9300 = 9'h140 == r_count_22_io_out ? io_r_320_b : _GEN_9299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9301 = 9'h141 == r_count_22_io_out ? io_r_321_b : _GEN_9300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9302 = 9'h142 == r_count_22_io_out ? io_r_322_b : _GEN_9301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9303 = 9'h143 == r_count_22_io_out ? io_r_323_b : _GEN_9302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9304 = 9'h144 == r_count_22_io_out ? io_r_324_b : _GEN_9303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9305 = 9'h145 == r_count_22_io_out ? io_r_325_b : _GEN_9304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9306 = 9'h146 == r_count_22_io_out ? io_r_326_b : _GEN_9305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9307 = 9'h147 == r_count_22_io_out ? io_r_327_b : _GEN_9306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9308 = 9'h148 == r_count_22_io_out ? io_r_328_b : _GEN_9307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9309 = 9'h149 == r_count_22_io_out ? io_r_329_b : _GEN_9308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9310 = 9'h14a == r_count_22_io_out ? io_r_330_b : _GEN_9309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9311 = 9'h14b == r_count_22_io_out ? io_r_331_b : _GEN_9310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9312 = 9'h14c == r_count_22_io_out ? io_r_332_b : _GEN_9311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9313 = 9'h14d == r_count_22_io_out ? io_r_333_b : _GEN_9312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9314 = 9'h14e == r_count_22_io_out ? io_r_334_b : _GEN_9313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9315 = 9'h14f == r_count_22_io_out ? io_r_335_b : _GEN_9314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9316 = 9'h150 == r_count_22_io_out ? io_r_336_b : _GEN_9315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9317 = 9'h151 == r_count_22_io_out ? io_r_337_b : _GEN_9316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9318 = 9'h152 == r_count_22_io_out ? io_r_338_b : _GEN_9317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9319 = 9'h153 == r_count_22_io_out ? io_r_339_b : _GEN_9318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9320 = 9'h154 == r_count_22_io_out ? io_r_340_b : _GEN_9319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9321 = 9'h155 == r_count_22_io_out ? io_r_341_b : _GEN_9320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9322 = 9'h156 == r_count_22_io_out ? io_r_342_b : _GEN_9321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9323 = 9'h157 == r_count_22_io_out ? io_r_343_b : _GEN_9322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9324 = 9'h158 == r_count_22_io_out ? io_r_344_b : _GEN_9323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9325 = 9'h159 == r_count_22_io_out ? io_r_345_b : _GEN_9324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9326 = 9'h15a == r_count_22_io_out ? io_r_346_b : _GEN_9325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9327 = 9'h15b == r_count_22_io_out ? io_r_347_b : _GEN_9326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9328 = 9'h15c == r_count_22_io_out ? io_r_348_b : _GEN_9327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9329 = 9'h15d == r_count_22_io_out ? io_r_349_b : _GEN_9328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9330 = 9'h15e == r_count_22_io_out ? io_r_350_b : _GEN_9329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9331 = 9'h15f == r_count_22_io_out ? io_r_351_b : _GEN_9330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9332 = 9'h160 == r_count_22_io_out ? io_r_352_b : _GEN_9331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9333 = 9'h161 == r_count_22_io_out ? io_r_353_b : _GEN_9332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9334 = 9'h162 == r_count_22_io_out ? io_r_354_b : _GEN_9333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9335 = 9'h163 == r_count_22_io_out ? io_r_355_b : _GEN_9334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9336 = 9'h164 == r_count_22_io_out ? io_r_356_b : _GEN_9335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9337 = 9'h165 == r_count_22_io_out ? io_r_357_b : _GEN_9336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9338 = 9'h166 == r_count_22_io_out ? io_r_358_b : _GEN_9337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9339 = 9'h167 == r_count_22_io_out ? io_r_359_b : _GEN_9338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9340 = 9'h168 == r_count_22_io_out ? io_r_360_b : _GEN_9339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9341 = 9'h169 == r_count_22_io_out ? io_r_361_b : _GEN_9340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9342 = 9'h16a == r_count_22_io_out ? io_r_362_b : _GEN_9341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9343 = 9'h16b == r_count_22_io_out ? io_r_363_b : _GEN_9342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9344 = 9'h16c == r_count_22_io_out ? io_r_364_b : _GEN_9343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9345 = 9'h16d == r_count_22_io_out ? io_r_365_b : _GEN_9344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9346 = 9'h16e == r_count_22_io_out ? io_r_366_b : _GEN_9345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9347 = 9'h16f == r_count_22_io_out ? io_r_367_b : _GEN_9346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9348 = 9'h170 == r_count_22_io_out ? io_r_368_b : _GEN_9347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9349 = 9'h171 == r_count_22_io_out ? io_r_369_b : _GEN_9348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9350 = 9'h172 == r_count_22_io_out ? io_r_370_b : _GEN_9349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9351 = 9'h173 == r_count_22_io_out ? io_r_371_b : _GEN_9350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9352 = 9'h174 == r_count_22_io_out ? io_r_372_b : _GEN_9351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9353 = 9'h175 == r_count_22_io_out ? io_r_373_b : _GEN_9352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9354 = 9'h176 == r_count_22_io_out ? io_r_374_b : _GEN_9353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9355 = 9'h177 == r_count_22_io_out ? io_r_375_b : _GEN_9354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9356 = 9'h178 == r_count_22_io_out ? io_r_376_b : _GEN_9355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9357 = 9'h179 == r_count_22_io_out ? io_r_377_b : _GEN_9356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9358 = 9'h17a == r_count_22_io_out ? io_r_378_b : _GEN_9357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9359 = 9'h17b == r_count_22_io_out ? io_r_379_b : _GEN_9358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9360 = 9'h17c == r_count_22_io_out ? io_r_380_b : _GEN_9359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9361 = 9'h17d == r_count_22_io_out ? io_r_381_b : _GEN_9360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9362 = 9'h17e == r_count_22_io_out ? io_r_382_b : _GEN_9361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9363 = 9'h17f == r_count_22_io_out ? io_r_383_b : _GEN_9362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9364 = 9'h180 == r_count_22_io_out ? io_r_384_b : _GEN_9363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9365 = 9'h181 == r_count_22_io_out ? io_r_385_b : _GEN_9364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9366 = 9'h182 == r_count_22_io_out ? io_r_386_b : _GEN_9365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9367 = 9'h183 == r_count_22_io_out ? io_r_387_b : _GEN_9366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9368 = 9'h184 == r_count_22_io_out ? io_r_388_b : _GEN_9367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9369 = 9'h185 == r_count_22_io_out ? io_r_389_b : _GEN_9368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9370 = 9'h186 == r_count_22_io_out ? io_r_390_b : _GEN_9369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9371 = 9'h187 == r_count_22_io_out ? io_r_391_b : _GEN_9370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9372 = 9'h188 == r_count_22_io_out ? io_r_392_b : _GEN_9371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9373 = 9'h189 == r_count_22_io_out ? io_r_393_b : _GEN_9372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9374 = 9'h18a == r_count_22_io_out ? io_r_394_b : _GEN_9373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9375 = 9'h18b == r_count_22_io_out ? io_r_395_b : _GEN_9374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9376 = 9'h18c == r_count_22_io_out ? io_r_396_b : _GEN_9375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9377 = 9'h18d == r_count_22_io_out ? io_r_397_b : _GEN_9376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9378 = 9'h18e == r_count_22_io_out ? io_r_398_b : _GEN_9377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9381 = 9'h1 == r_count_23_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9382 = 9'h2 == r_count_23_io_out ? io_r_2_b : _GEN_9381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9383 = 9'h3 == r_count_23_io_out ? io_r_3_b : _GEN_9382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9384 = 9'h4 == r_count_23_io_out ? io_r_4_b : _GEN_9383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9385 = 9'h5 == r_count_23_io_out ? io_r_5_b : _GEN_9384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9386 = 9'h6 == r_count_23_io_out ? io_r_6_b : _GEN_9385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9387 = 9'h7 == r_count_23_io_out ? io_r_7_b : _GEN_9386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9388 = 9'h8 == r_count_23_io_out ? io_r_8_b : _GEN_9387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9389 = 9'h9 == r_count_23_io_out ? io_r_9_b : _GEN_9388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9390 = 9'ha == r_count_23_io_out ? io_r_10_b : _GEN_9389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9391 = 9'hb == r_count_23_io_out ? io_r_11_b : _GEN_9390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9392 = 9'hc == r_count_23_io_out ? io_r_12_b : _GEN_9391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9393 = 9'hd == r_count_23_io_out ? io_r_13_b : _GEN_9392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9394 = 9'he == r_count_23_io_out ? io_r_14_b : _GEN_9393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9395 = 9'hf == r_count_23_io_out ? io_r_15_b : _GEN_9394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9396 = 9'h10 == r_count_23_io_out ? io_r_16_b : _GEN_9395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9397 = 9'h11 == r_count_23_io_out ? io_r_17_b : _GEN_9396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9398 = 9'h12 == r_count_23_io_out ? io_r_18_b : _GEN_9397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9399 = 9'h13 == r_count_23_io_out ? io_r_19_b : _GEN_9398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9400 = 9'h14 == r_count_23_io_out ? io_r_20_b : _GEN_9399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9401 = 9'h15 == r_count_23_io_out ? io_r_21_b : _GEN_9400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9402 = 9'h16 == r_count_23_io_out ? io_r_22_b : _GEN_9401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9403 = 9'h17 == r_count_23_io_out ? io_r_23_b : _GEN_9402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9404 = 9'h18 == r_count_23_io_out ? io_r_24_b : _GEN_9403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9405 = 9'h19 == r_count_23_io_out ? io_r_25_b : _GEN_9404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9406 = 9'h1a == r_count_23_io_out ? io_r_26_b : _GEN_9405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9407 = 9'h1b == r_count_23_io_out ? io_r_27_b : _GEN_9406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9408 = 9'h1c == r_count_23_io_out ? io_r_28_b : _GEN_9407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9409 = 9'h1d == r_count_23_io_out ? io_r_29_b : _GEN_9408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9410 = 9'h1e == r_count_23_io_out ? io_r_30_b : _GEN_9409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9411 = 9'h1f == r_count_23_io_out ? io_r_31_b : _GEN_9410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9412 = 9'h20 == r_count_23_io_out ? io_r_32_b : _GEN_9411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9413 = 9'h21 == r_count_23_io_out ? io_r_33_b : _GEN_9412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9414 = 9'h22 == r_count_23_io_out ? io_r_34_b : _GEN_9413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9415 = 9'h23 == r_count_23_io_out ? io_r_35_b : _GEN_9414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9416 = 9'h24 == r_count_23_io_out ? io_r_36_b : _GEN_9415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9417 = 9'h25 == r_count_23_io_out ? io_r_37_b : _GEN_9416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9418 = 9'h26 == r_count_23_io_out ? io_r_38_b : _GEN_9417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9419 = 9'h27 == r_count_23_io_out ? io_r_39_b : _GEN_9418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9420 = 9'h28 == r_count_23_io_out ? io_r_40_b : _GEN_9419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9421 = 9'h29 == r_count_23_io_out ? io_r_41_b : _GEN_9420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9422 = 9'h2a == r_count_23_io_out ? io_r_42_b : _GEN_9421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9423 = 9'h2b == r_count_23_io_out ? io_r_43_b : _GEN_9422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9424 = 9'h2c == r_count_23_io_out ? io_r_44_b : _GEN_9423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9425 = 9'h2d == r_count_23_io_out ? io_r_45_b : _GEN_9424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9426 = 9'h2e == r_count_23_io_out ? io_r_46_b : _GEN_9425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9427 = 9'h2f == r_count_23_io_out ? io_r_47_b : _GEN_9426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9428 = 9'h30 == r_count_23_io_out ? io_r_48_b : _GEN_9427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9429 = 9'h31 == r_count_23_io_out ? io_r_49_b : _GEN_9428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9430 = 9'h32 == r_count_23_io_out ? io_r_50_b : _GEN_9429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9431 = 9'h33 == r_count_23_io_out ? io_r_51_b : _GEN_9430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9432 = 9'h34 == r_count_23_io_out ? io_r_52_b : _GEN_9431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9433 = 9'h35 == r_count_23_io_out ? io_r_53_b : _GEN_9432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9434 = 9'h36 == r_count_23_io_out ? io_r_54_b : _GEN_9433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9435 = 9'h37 == r_count_23_io_out ? io_r_55_b : _GEN_9434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9436 = 9'h38 == r_count_23_io_out ? io_r_56_b : _GEN_9435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9437 = 9'h39 == r_count_23_io_out ? io_r_57_b : _GEN_9436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9438 = 9'h3a == r_count_23_io_out ? io_r_58_b : _GEN_9437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9439 = 9'h3b == r_count_23_io_out ? io_r_59_b : _GEN_9438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9440 = 9'h3c == r_count_23_io_out ? io_r_60_b : _GEN_9439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9441 = 9'h3d == r_count_23_io_out ? io_r_61_b : _GEN_9440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9442 = 9'h3e == r_count_23_io_out ? io_r_62_b : _GEN_9441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9443 = 9'h3f == r_count_23_io_out ? io_r_63_b : _GEN_9442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9444 = 9'h40 == r_count_23_io_out ? io_r_64_b : _GEN_9443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9445 = 9'h41 == r_count_23_io_out ? io_r_65_b : _GEN_9444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9446 = 9'h42 == r_count_23_io_out ? io_r_66_b : _GEN_9445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9447 = 9'h43 == r_count_23_io_out ? io_r_67_b : _GEN_9446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9448 = 9'h44 == r_count_23_io_out ? io_r_68_b : _GEN_9447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9449 = 9'h45 == r_count_23_io_out ? io_r_69_b : _GEN_9448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9450 = 9'h46 == r_count_23_io_out ? io_r_70_b : _GEN_9449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9451 = 9'h47 == r_count_23_io_out ? io_r_71_b : _GEN_9450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9452 = 9'h48 == r_count_23_io_out ? io_r_72_b : _GEN_9451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9453 = 9'h49 == r_count_23_io_out ? io_r_73_b : _GEN_9452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9454 = 9'h4a == r_count_23_io_out ? io_r_74_b : _GEN_9453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9455 = 9'h4b == r_count_23_io_out ? io_r_75_b : _GEN_9454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9456 = 9'h4c == r_count_23_io_out ? io_r_76_b : _GEN_9455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9457 = 9'h4d == r_count_23_io_out ? io_r_77_b : _GEN_9456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9458 = 9'h4e == r_count_23_io_out ? io_r_78_b : _GEN_9457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9459 = 9'h4f == r_count_23_io_out ? io_r_79_b : _GEN_9458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9460 = 9'h50 == r_count_23_io_out ? io_r_80_b : _GEN_9459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9461 = 9'h51 == r_count_23_io_out ? io_r_81_b : _GEN_9460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9462 = 9'h52 == r_count_23_io_out ? io_r_82_b : _GEN_9461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9463 = 9'h53 == r_count_23_io_out ? io_r_83_b : _GEN_9462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9464 = 9'h54 == r_count_23_io_out ? io_r_84_b : _GEN_9463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9465 = 9'h55 == r_count_23_io_out ? io_r_85_b : _GEN_9464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9466 = 9'h56 == r_count_23_io_out ? io_r_86_b : _GEN_9465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9467 = 9'h57 == r_count_23_io_out ? io_r_87_b : _GEN_9466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9468 = 9'h58 == r_count_23_io_out ? io_r_88_b : _GEN_9467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9469 = 9'h59 == r_count_23_io_out ? io_r_89_b : _GEN_9468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9470 = 9'h5a == r_count_23_io_out ? io_r_90_b : _GEN_9469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9471 = 9'h5b == r_count_23_io_out ? io_r_91_b : _GEN_9470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9472 = 9'h5c == r_count_23_io_out ? io_r_92_b : _GEN_9471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9473 = 9'h5d == r_count_23_io_out ? io_r_93_b : _GEN_9472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9474 = 9'h5e == r_count_23_io_out ? io_r_94_b : _GEN_9473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9475 = 9'h5f == r_count_23_io_out ? io_r_95_b : _GEN_9474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9476 = 9'h60 == r_count_23_io_out ? io_r_96_b : _GEN_9475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9477 = 9'h61 == r_count_23_io_out ? io_r_97_b : _GEN_9476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9478 = 9'h62 == r_count_23_io_out ? io_r_98_b : _GEN_9477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9479 = 9'h63 == r_count_23_io_out ? io_r_99_b : _GEN_9478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9480 = 9'h64 == r_count_23_io_out ? io_r_100_b : _GEN_9479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9481 = 9'h65 == r_count_23_io_out ? io_r_101_b : _GEN_9480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9482 = 9'h66 == r_count_23_io_out ? io_r_102_b : _GEN_9481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9483 = 9'h67 == r_count_23_io_out ? io_r_103_b : _GEN_9482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9484 = 9'h68 == r_count_23_io_out ? io_r_104_b : _GEN_9483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9485 = 9'h69 == r_count_23_io_out ? io_r_105_b : _GEN_9484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9486 = 9'h6a == r_count_23_io_out ? io_r_106_b : _GEN_9485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9487 = 9'h6b == r_count_23_io_out ? io_r_107_b : _GEN_9486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9488 = 9'h6c == r_count_23_io_out ? io_r_108_b : _GEN_9487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9489 = 9'h6d == r_count_23_io_out ? io_r_109_b : _GEN_9488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9490 = 9'h6e == r_count_23_io_out ? io_r_110_b : _GEN_9489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9491 = 9'h6f == r_count_23_io_out ? io_r_111_b : _GEN_9490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9492 = 9'h70 == r_count_23_io_out ? io_r_112_b : _GEN_9491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9493 = 9'h71 == r_count_23_io_out ? io_r_113_b : _GEN_9492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9494 = 9'h72 == r_count_23_io_out ? io_r_114_b : _GEN_9493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9495 = 9'h73 == r_count_23_io_out ? io_r_115_b : _GEN_9494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9496 = 9'h74 == r_count_23_io_out ? io_r_116_b : _GEN_9495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9497 = 9'h75 == r_count_23_io_out ? io_r_117_b : _GEN_9496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9498 = 9'h76 == r_count_23_io_out ? io_r_118_b : _GEN_9497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9499 = 9'h77 == r_count_23_io_out ? io_r_119_b : _GEN_9498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9500 = 9'h78 == r_count_23_io_out ? io_r_120_b : _GEN_9499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9501 = 9'h79 == r_count_23_io_out ? io_r_121_b : _GEN_9500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9502 = 9'h7a == r_count_23_io_out ? io_r_122_b : _GEN_9501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9503 = 9'h7b == r_count_23_io_out ? io_r_123_b : _GEN_9502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9504 = 9'h7c == r_count_23_io_out ? io_r_124_b : _GEN_9503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9505 = 9'h7d == r_count_23_io_out ? io_r_125_b : _GEN_9504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9506 = 9'h7e == r_count_23_io_out ? io_r_126_b : _GEN_9505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9507 = 9'h7f == r_count_23_io_out ? io_r_127_b : _GEN_9506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9508 = 9'h80 == r_count_23_io_out ? io_r_128_b : _GEN_9507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9509 = 9'h81 == r_count_23_io_out ? io_r_129_b : _GEN_9508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9510 = 9'h82 == r_count_23_io_out ? io_r_130_b : _GEN_9509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9511 = 9'h83 == r_count_23_io_out ? io_r_131_b : _GEN_9510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9512 = 9'h84 == r_count_23_io_out ? io_r_132_b : _GEN_9511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9513 = 9'h85 == r_count_23_io_out ? io_r_133_b : _GEN_9512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9514 = 9'h86 == r_count_23_io_out ? io_r_134_b : _GEN_9513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9515 = 9'h87 == r_count_23_io_out ? io_r_135_b : _GEN_9514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9516 = 9'h88 == r_count_23_io_out ? io_r_136_b : _GEN_9515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9517 = 9'h89 == r_count_23_io_out ? io_r_137_b : _GEN_9516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9518 = 9'h8a == r_count_23_io_out ? io_r_138_b : _GEN_9517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9519 = 9'h8b == r_count_23_io_out ? io_r_139_b : _GEN_9518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9520 = 9'h8c == r_count_23_io_out ? io_r_140_b : _GEN_9519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9521 = 9'h8d == r_count_23_io_out ? io_r_141_b : _GEN_9520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9522 = 9'h8e == r_count_23_io_out ? io_r_142_b : _GEN_9521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9523 = 9'h8f == r_count_23_io_out ? io_r_143_b : _GEN_9522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9524 = 9'h90 == r_count_23_io_out ? io_r_144_b : _GEN_9523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9525 = 9'h91 == r_count_23_io_out ? io_r_145_b : _GEN_9524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9526 = 9'h92 == r_count_23_io_out ? io_r_146_b : _GEN_9525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9527 = 9'h93 == r_count_23_io_out ? io_r_147_b : _GEN_9526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9528 = 9'h94 == r_count_23_io_out ? io_r_148_b : _GEN_9527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9529 = 9'h95 == r_count_23_io_out ? io_r_149_b : _GEN_9528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9530 = 9'h96 == r_count_23_io_out ? io_r_150_b : _GEN_9529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9531 = 9'h97 == r_count_23_io_out ? io_r_151_b : _GEN_9530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9532 = 9'h98 == r_count_23_io_out ? io_r_152_b : _GEN_9531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9533 = 9'h99 == r_count_23_io_out ? io_r_153_b : _GEN_9532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9534 = 9'h9a == r_count_23_io_out ? io_r_154_b : _GEN_9533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9535 = 9'h9b == r_count_23_io_out ? io_r_155_b : _GEN_9534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9536 = 9'h9c == r_count_23_io_out ? io_r_156_b : _GEN_9535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9537 = 9'h9d == r_count_23_io_out ? io_r_157_b : _GEN_9536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9538 = 9'h9e == r_count_23_io_out ? io_r_158_b : _GEN_9537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9539 = 9'h9f == r_count_23_io_out ? io_r_159_b : _GEN_9538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9540 = 9'ha0 == r_count_23_io_out ? io_r_160_b : _GEN_9539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9541 = 9'ha1 == r_count_23_io_out ? io_r_161_b : _GEN_9540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9542 = 9'ha2 == r_count_23_io_out ? io_r_162_b : _GEN_9541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9543 = 9'ha3 == r_count_23_io_out ? io_r_163_b : _GEN_9542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9544 = 9'ha4 == r_count_23_io_out ? io_r_164_b : _GEN_9543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9545 = 9'ha5 == r_count_23_io_out ? io_r_165_b : _GEN_9544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9546 = 9'ha6 == r_count_23_io_out ? io_r_166_b : _GEN_9545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9547 = 9'ha7 == r_count_23_io_out ? io_r_167_b : _GEN_9546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9548 = 9'ha8 == r_count_23_io_out ? io_r_168_b : _GEN_9547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9549 = 9'ha9 == r_count_23_io_out ? io_r_169_b : _GEN_9548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9550 = 9'haa == r_count_23_io_out ? io_r_170_b : _GEN_9549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9551 = 9'hab == r_count_23_io_out ? io_r_171_b : _GEN_9550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9552 = 9'hac == r_count_23_io_out ? io_r_172_b : _GEN_9551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9553 = 9'had == r_count_23_io_out ? io_r_173_b : _GEN_9552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9554 = 9'hae == r_count_23_io_out ? io_r_174_b : _GEN_9553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9555 = 9'haf == r_count_23_io_out ? io_r_175_b : _GEN_9554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9556 = 9'hb0 == r_count_23_io_out ? io_r_176_b : _GEN_9555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9557 = 9'hb1 == r_count_23_io_out ? io_r_177_b : _GEN_9556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9558 = 9'hb2 == r_count_23_io_out ? io_r_178_b : _GEN_9557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9559 = 9'hb3 == r_count_23_io_out ? io_r_179_b : _GEN_9558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9560 = 9'hb4 == r_count_23_io_out ? io_r_180_b : _GEN_9559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9561 = 9'hb5 == r_count_23_io_out ? io_r_181_b : _GEN_9560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9562 = 9'hb6 == r_count_23_io_out ? io_r_182_b : _GEN_9561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9563 = 9'hb7 == r_count_23_io_out ? io_r_183_b : _GEN_9562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9564 = 9'hb8 == r_count_23_io_out ? io_r_184_b : _GEN_9563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9565 = 9'hb9 == r_count_23_io_out ? io_r_185_b : _GEN_9564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9566 = 9'hba == r_count_23_io_out ? io_r_186_b : _GEN_9565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9567 = 9'hbb == r_count_23_io_out ? io_r_187_b : _GEN_9566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9568 = 9'hbc == r_count_23_io_out ? io_r_188_b : _GEN_9567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9569 = 9'hbd == r_count_23_io_out ? io_r_189_b : _GEN_9568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9570 = 9'hbe == r_count_23_io_out ? io_r_190_b : _GEN_9569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9571 = 9'hbf == r_count_23_io_out ? io_r_191_b : _GEN_9570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9572 = 9'hc0 == r_count_23_io_out ? io_r_192_b : _GEN_9571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9573 = 9'hc1 == r_count_23_io_out ? io_r_193_b : _GEN_9572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9574 = 9'hc2 == r_count_23_io_out ? io_r_194_b : _GEN_9573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9575 = 9'hc3 == r_count_23_io_out ? io_r_195_b : _GEN_9574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9576 = 9'hc4 == r_count_23_io_out ? io_r_196_b : _GEN_9575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9577 = 9'hc5 == r_count_23_io_out ? io_r_197_b : _GEN_9576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9578 = 9'hc6 == r_count_23_io_out ? io_r_198_b : _GEN_9577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9579 = 9'hc7 == r_count_23_io_out ? io_r_199_b : _GEN_9578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9580 = 9'hc8 == r_count_23_io_out ? io_r_200_b : _GEN_9579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9581 = 9'hc9 == r_count_23_io_out ? io_r_201_b : _GEN_9580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9582 = 9'hca == r_count_23_io_out ? io_r_202_b : _GEN_9581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9583 = 9'hcb == r_count_23_io_out ? io_r_203_b : _GEN_9582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9584 = 9'hcc == r_count_23_io_out ? io_r_204_b : _GEN_9583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9585 = 9'hcd == r_count_23_io_out ? io_r_205_b : _GEN_9584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9586 = 9'hce == r_count_23_io_out ? io_r_206_b : _GEN_9585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9587 = 9'hcf == r_count_23_io_out ? io_r_207_b : _GEN_9586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9588 = 9'hd0 == r_count_23_io_out ? io_r_208_b : _GEN_9587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9589 = 9'hd1 == r_count_23_io_out ? io_r_209_b : _GEN_9588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9590 = 9'hd2 == r_count_23_io_out ? io_r_210_b : _GEN_9589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9591 = 9'hd3 == r_count_23_io_out ? io_r_211_b : _GEN_9590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9592 = 9'hd4 == r_count_23_io_out ? io_r_212_b : _GEN_9591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9593 = 9'hd5 == r_count_23_io_out ? io_r_213_b : _GEN_9592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9594 = 9'hd6 == r_count_23_io_out ? io_r_214_b : _GEN_9593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9595 = 9'hd7 == r_count_23_io_out ? io_r_215_b : _GEN_9594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9596 = 9'hd8 == r_count_23_io_out ? io_r_216_b : _GEN_9595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9597 = 9'hd9 == r_count_23_io_out ? io_r_217_b : _GEN_9596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9598 = 9'hda == r_count_23_io_out ? io_r_218_b : _GEN_9597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9599 = 9'hdb == r_count_23_io_out ? io_r_219_b : _GEN_9598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9600 = 9'hdc == r_count_23_io_out ? io_r_220_b : _GEN_9599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9601 = 9'hdd == r_count_23_io_out ? io_r_221_b : _GEN_9600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9602 = 9'hde == r_count_23_io_out ? io_r_222_b : _GEN_9601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9603 = 9'hdf == r_count_23_io_out ? io_r_223_b : _GEN_9602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9604 = 9'he0 == r_count_23_io_out ? io_r_224_b : _GEN_9603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9605 = 9'he1 == r_count_23_io_out ? io_r_225_b : _GEN_9604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9606 = 9'he2 == r_count_23_io_out ? io_r_226_b : _GEN_9605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9607 = 9'he3 == r_count_23_io_out ? io_r_227_b : _GEN_9606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9608 = 9'he4 == r_count_23_io_out ? io_r_228_b : _GEN_9607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9609 = 9'he5 == r_count_23_io_out ? io_r_229_b : _GEN_9608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9610 = 9'he6 == r_count_23_io_out ? io_r_230_b : _GEN_9609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9611 = 9'he7 == r_count_23_io_out ? io_r_231_b : _GEN_9610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9612 = 9'he8 == r_count_23_io_out ? io_r_232_b : _GEN_9611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9613 = 9'he9 == r_count_23_io_out ? io_r_233_b : _GEN_9612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9614 = 9'hea == r_count_23_io_out ? io_r_234_b : _GEN_9613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9615 = 9'heb == r_count_23_io_out ? io_r_235_b : _GEN_9614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9616 = 9'hec == r_count_23_io_out ? io_r_236_b : _GEN_9615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9617 = 9'hed == r_count_23_io_out ? io_r_237_b : _GEN_9616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9618 = 9'hee == r_count_23_io_out ? io_r_238_b : _GEN_9617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9619 = 9'hef == r_count_23_io_out ? io_r_239_b : _GEN_9618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9620 = 9'hf0 == r_count_23_io_out ? io_r_240_b : _GEN_9619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9621 = 9'hf1 == r_count_23_io_out ? io_r_241_b : _GEN_9620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9622 = 9'hf2 == r_count_23_io_out ? io_r_242_b : _GEN_9621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9623 = 9'hf3 == r_count_23_io_out ? io_r_243_b : _GEN_9622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9624 = 9'hf4 == r_count_23_io_out ? io_r_244_b : _GEN_9623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9625 = 9'hf5 == r_count_23_io_out ? io_r_245_b : _GEN_9624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9626 = 9'hf6 == r_count_23_io_out ? io_r_246_b : _GEN_9625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9627 = 9'hf7 == r_count_23_io_out ? io_r_247_b : _GEN_9626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9628 = 9'hf8 == r_count_23_io_out ? io_r_248_b : _GEN_9627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9629 = 9'hf9 == r_count_23_io_out ? io_r_249_b : _GEN_9628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9630 = 9'hfa == r_count_23_io_out ? io_r_250_b : _GEN_9629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9631 = 9'hfb == r_count_23_io_out ? io_r_251_b : _GEN_9630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9632 = 9'hfc == r_count_23_io_out ? io_r_252_b : _GEN_9631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9633 = 9'hfd == r_count_23_io_out ? io_r_253_b : _GEN_9632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9634 = 9'hfe == r_count_23_io_out ? io_r_254_b : _GEN_9633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9635 = 9'hff == r_count_23_io_out ? io_r_255_b : _GEN_9634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9636 = 9'h100 == r_count_23_io_out ? io_r_256_b : _GEN_9635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9637 = 9'h101 == r_count_23_io_out ? io_r_257_b : _GEN_9636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9638 = 9'h102 == r_count_23_io_out ? io_r_258_b : _GEN_9637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9639 = 9'h103 == r_count_23_io_out ? io_r_259_b : _GEN_9638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9640 = 9'h104 == r_count_23_io_out ? io_r_260_b : _GEN_9639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9641 = 9'h105 == r_count_23_io_out ? io_r_261_b : _GEN_9640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9642 = 9'h106 == r_count_23_io_out ? io_r_262_b : _GEN_9641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9643 = 9'h107 == r_count_23_io_out ? io_r_263_b : _GEN_9642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9644 = 9'h108 == r_count_23_io_out ? io_r_264_b : _GEN_9643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9645 = 9'h109 == r_count_23_io_out ? io_r_265_b : _GEN_9644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9646 = 9'h10a == r_count_23_io_out ? io_r_266_b : _GEN_9645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9647 = 9'h10b == r_count_23_io_out ? io_r_267_b : _GEN_9646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9648 = 9'h10c == r_count_23_io_out ? io_r_268_b : _GEN_9647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9649 = 9'h10d == r_count_23_io_out ? io_r_269_b : _GEN_9648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9650 = 9'h10e == r_count_23_io_out ? io_r_270_b : _GEN_9649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9651 = 9'h10f == r_count_23_io_out ? io_r_271_b : _GEN_9650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9652 = 9'h110 == r_count_23_io_out ? io_r_272_b : _GEN_9651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9653 = 9'h111 == r_count_23_io_out ? io_r_273_b : _GEN_9652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9654 = 9'h112 == r_count_23_io_out ? io_r_274_b : _GEN_9653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9655 = 9'h113 == r_count_23_io_out ? io_r_275_b : _GEN_9654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9656 = 9'h114 == r_count_23_io_out ? io_r_276_b : _GEN_9655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9657 = 9'h115 == r_count_23_io_out ? io_r_277_b : _GEN_9656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9658 = 9'h116 == r_count_23_io_out ? io_r_278_b : _GEN_9657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9659 = 9'h117 == r_count_23_io_out ? io_r_279_b : _GEN_9658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9660 = 9'h118 == r_count_23_io_out ? io_r_280_b : _GEN_9659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9661 = 9'h119 == r_count_23_io_out ? io_r_281_b : _GEN_9660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9662 = 9'h11a == r_count_23_io_out ? io_r_282_b : _GEN_9661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9663 = 9'h11b == r_count_23_io_out ? io_r_283_b : _GEN_9662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9664 = 9'h11c == r_count_23_io_out ? io_r_284_b : _GEN_9663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9665 = 9'h11d == r_count_23_io_out ? io_r_285_b : _GEN_9664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9666 = 9'h11e == r_count_23_io_out ? io_r_286_b : _GEN_9665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9667 = 9'h11f == r_count_23_io_out ? io_r_287_b : _GEN_9666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9668 = 9'h120 == r_count_23_io_out ? io_r_288_b : _GEN_9667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9669 = 9'h121 == r_count_23_io_out ? io_r_289_b : _GEN_9668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9670 = 9'h122 == r_count_23_io_out ? io_r_290_b : _GEN_9669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9671 = 9'h123 == r_count_23_io_out ? io_r_291_b : _GEN_9670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9672 = 9'h124 == r_count_23_io_out ? io_r_292_b : _GEN_9671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9673 = 9'h125 == r_count_23_io_out ? io_r_293_b : _GEN_9672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9674 = 9'h126 == r_count_23_io_out ? io_r_294_b : _GEN_9673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9675 = 9'h127 == r_count_23_io_out ? io_r_295_b : _GEN_9674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9676 = 9'h128 == r_count_23_io_out ? io_r_296_b : _GEN_9675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9677 = 9'h129 == r_count_23_io_out ? io_r_297_b : _GEN_9676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9678 = 9'h12a == r_count_23_io_out ? io_r_298_b : _GEN_9677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9679 = 9'h12b == r_count_23_io_out ? io_r_299_b : _GEN_9678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9680 = 9'h12c == r_count_23_io_out ? io_r_300_b : _GEN_9679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9681 = 9'h12d == r_count_23_io_out ? io_r_301_b : _GEN_9680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9682 = 9'h12e == r_count_23_io_out ? io_r_302_b : _GEN_9681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9683 = 9'h12f == r_count_23_io_out ? io_r_303_b : _GEN_9682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9684 = 9'h130 == r_count_23_io_out ? io_r_304_b : _GEN_9683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9685 = 9'h131 == r_count_23_io_out ? io_r_305_b : _GEN_9684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9686 = 9'h132 == r_count_23_io_out ? io_r_306_b : _GEN_9685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9687 = 9'h133 == r_count_23_io_out ? io_r_307_b : _GEN_9686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9688 = 9'h134 == r_count_23_io_out ? io_r_308_b : _GEN_9687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9689 = 9'h135 == r_count_23_io_out ? io_r_309_b : _GEN_9688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9690 = 9'h136 == r_count_23_io_out ? io_r_310_b : _GEN_9689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9691 = 9'h137 == r_count_23_io_out ? io_r_311_b : _GEN_9690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9692 = 9'h138 == r_count_23_io_out ? io_r_312_b : _GEN_9691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9693 = 9'h139 == r_count_23_io_out ? io_r_313_b : _GEN_9692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9694 = 9'h13a == r_count_23_io_out ? io_r_314_b : _GEN_9693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9695 = 9'h13b == r_count_23_io_out ? io_r_315_b : _GEN_9694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9696 = 9'h13c == r_count_23_io_out ? io_r_316_b : _GEN_9695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9697 = 9'h13d == r_count_23_io_out ? io_r_317_b : _GEN_9696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9698 = 9'h13e == r_count_23_io_out ? io_r_318_b : _GEN_9697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9699 = 9'h13f == r_count_23_io_out ? io_r_319_b : _GEN_9698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9700 = 9'h140 == r_count_23_io_out ? io_r_320_b : _GEN_9699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9701 = 9'h141 == r_count_23_io_out ? io_r_321_b : _GEN_9700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9702 = 9'h142 == r_count_23_io_out ? io_r_322_b : _GEN_9701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9703 = 9'h143 == r_count_23_io_out ? io_r_323_b : _GEN_9702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9704 = 9'h144 == r_count_23_io_out ? io_r_324_b : _GEN_9703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9705 = 9'h145 == r_count_23_io_out ? io_r_325_b : _GEN_9704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9706 = 9'h146 == r_count_23_io_out ? io_r_326_b : _GEN_9705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9707 = 9'h147 == r_count_23_io_out ? io_r_327_b : _GEN_9706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9708 = 9'h148 == r_count_23_io_out ? io_r_328_b : _GEN_9707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9709 = 9'h149 == r_count_23_io_out ? io_r_329_b : _GEN_9708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9710 = 9'h14a == r_count_23_io_out ? io_r_330_b : _GEN_9709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9711 = 9'h14b == r_count_23_io_out ? io_r_331_b : _GEN_9710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9712 = 9'h14c == r_count_23_io_out ? io_r_332_b : _GEN_9711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9713 = 9'h14d == r_count_23_io_out ? io_r_333_b : _GEN_9712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9714 = 9'h14e == r_count_23_io_out ? io_r_334_b : _GEN_9713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9715 = 9'h14f == r_count_23_io_out ? io_r_335_b : _GEN_9714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9716 = 9'h150 == r_count_23_io_out ? io_r_336_b : _GEN_9715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9717 = 9'h151 == r_count_23_io_out ? io_r_337_b : _GEN_9716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9718 = 9'h152 == r_count_23_io_out ? io_r_338_b : _GEN_9717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9719 = 9'h153 == r_count_23_io_out ? io_r_339_b : _GEN_9718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9720 = 9'h154 == r_count_23_io_out ? io_r_340_b : _GEN_9719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9721 = 9'h155 == r_count_23_io_out ? io_r_341_b : _GEN_9720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9722 = 9'h156 == r_count_23_io_out ? io_r_342_b : _GEN_9721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9723 = 9'h157 == r_count_23_io_out ? io_r_343_b : _GEN_9722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9724 = 9'h158 == r_count_23_io_out ? io_r_344_b : _GEN_9723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9725 = 9'h159 == r_count_23_io_out ? io_r_345_b : _GEN_9724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9726 = 9'h15a == r_count_23_io_out ? io_r_346_b : _GEN_9725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9727 = 9'h15b == r_count_23_io_out ? io_r_347_b : _GEN_9726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9728 = 9'h15c == r_count_23_io_out ? io_r_348_b : _GEN_9727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9729 = 9'h15d == r_count_23_io_out ? io_r_349_b : _GEN_9728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9730 = 9'h15e == r_count_23_io_out ? io_r_350_b : _GEN_9729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9731 = 9'h15f == r_count_23_io_out ? io_r_351_b : _GEN_9730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9732 = 9'h160 == r_count_23_io_out ? io_r_352_b : _GEN_9731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9733 = 9'h161 == r_count_23_io_out ? io_r_353_b : _GEN_9732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9734 = 9'h162 == r_count_23_io_out ? io_r_354_b : _GEN_9733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9735 = 9'h163 == r_count_23_io_out ? io_r_355_b : _GEN_9734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9736 = 9'h164 == r_count_23_io_out ? io_r_356_b : _GEN_9735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9737 = 9'h165 == r_count_23_io_out ? io_r_357_b : _GEN_9736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9738 = 9'h166 == r_count_23_io_out ? io_r_358_b : _GEN_9737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9739 = 9'h167 == r_count_23_io_out ? io_r_359_b : _GEN_9738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9740 = 9'h168 == r_count_23_io_out ? io_r_360_b : _GEN_9739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9741 = 9'h169 == r_count_23_io_out ? io_r_361_b : _GEN_9740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9742 = 9'h16a == r_count_23_io_out ? io_r_362_b : _GEN_9741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9743 = 9'h16b == r_count_23_io_out ? io_r_363_b : _GEN_9742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9744 = 9'h16c == r_count_23_io_out ? io_r_364_b : _GEN_9743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9745 = 9'h16d == r_count_23_io_out ? io_r_365_b : _GEN_9744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9746 = 9'h16e == r_count_23_io_out ? io_r_366_b : _GEN_9745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9747 = 9'h16f == r_count_23_io_out ? io_r_367_b : _GEN_9746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9748 = 9'h170 == r_count_23_io_out ? io_r_368_b : _GEN_9747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9749 = 9'h171 == r_count_23_io_out ? io_r_369_b : _GEN_9748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9750 = 9'h172 == r_count_23_io_out ? io_r_370_b : _GEN_9749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9751 = 9'h173 == r_count_23_io_out ? io_r_371_b : _GEN_9750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9752 = 9'h174 == r_count_23_io_out ? io_r_372_b : _GEN_9751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9753 = 9'h175 == r_count_23_io_out ? io_r_373_b : _GEN_9752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9754 = 9'h176 == r_count_23_io_out ? io_r_374_b : _GEN_9753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9755 = 9'h177 == r_count_23_io_out ? io_r_375_b : _GEN_9754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9756 = 9'h178 == r_count_23_io_out ? io_r_376_b : _GEN_9755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9757 = 9'h179 == r_count_23_io_out ? io_r_377_b : _GEN_9756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9758 = 9'h17a == r_count_23_io_out ? io_r_378_b : _GEN_9757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9759 = 9'h17b == r_count_23_io_out ? io_r_379_b : _GEN_9758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9760 = 9'h17c == r_count_23_io_out ? io_r_380_b : _GEN_9759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9761 = 9'h17d == r_count_23_io_out ? io_r_381_b : _GEN_9760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9762 = 9'h17e == r_count_23_io_out ? io_r_382_b : _GEN_9761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9763 = 9'h17f == r_count_23_io_out ? io_r_383_b : _GEN_9762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9764 = 9'h180 == r_count_23_io_out ? io_r_384_b : _GEN_9763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9765 = 9'h181 == r_count_23_io_out ? io_r_385_b : _GEN_9764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9766 = 9'h182 == r_count_23_io_out ? io_r_386_b : _GEN_9765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9767 = 9'h183 == r_count_23_io_out ? io_r_387_b : _GEN_9766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9768 = 9'h184 == r_count_23_io_out ? io_r_388_b : _GEN_9767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9769 = 9'h185 == r_count_23_io_out ? io_r_389_b : _GEN_9768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9770 = 9'h186 == r_count_23_io_out ? io_r_390_b : _GEN_9769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9771 = 9'h187 == r_count_23_io_out ? io_r_391_b : _GEN_9770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9772 = 9'h188 == r_count_23_io_out ? io_r_392_b : _GEN_9771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9773 = 9'h189 == r_count_23_io_out ? io_r_393_b : _GEN_9772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9774 = 9'h18a == r_count_23_io_out ? io_r_394_b : _GEN_9773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9775 = 9'h18b == r_count_23_io_out ? io_r_395_b : _GEN_9774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9776 = 9'h18c == r_count_23_io_out ? io_r_396_b : _GEN_9775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9777 = 9'h18d == r_count_23_io_out ? io_r_397_b : _GEN_9776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9778 = 9'h18e == r_count_23_io_out ? io_r_398_b : _GEN_9777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9781 = 9'h1 == r_count_24_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9782 = 9'h2 == r_count_24_io_out ? io_r_2_b : _GEN_9781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9783 = 9'h3 == r_count_24_io_out ? io_r_3_b : _GEN_9782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9784 = 9'h4 == r_count_24_io_out ? io_r_4_b : _GEN_9783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9785 = 9'h5 == r_count_24_io_out ? io_r_5_b : _GEN_9784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9786 = 9'h6 == r_count_24_io_out ? io_r_6_b : _GEN_9785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9787 = 9'h7 == r_count_24_io_out ? io_r_7_b : _GEN_9786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9788 = 9'h8 == r_count_24_io_out ? io_r_8_b : _GEN_9787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9789 = 9'h9 == r_count_24_io_out ? io_r_9_b : _GEN_9788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9790 = 9'ha == r_count_24_io_out ? io_r_10_b : _GEN_9789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9791 = 9'hb == r_count_24_io_out ? io_r_11_b : _GEN_9790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9792 = 9'hc == r_count_24_io_out ? io_r_12_b : _GEN_9791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9793 = 9'hd == r_count_24_io_out ? io_r_13_b : _GEN_9792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9794 = 9'he == r_count_24_io_out ? io_r_14_b : _GEN_9793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9795 = 9'hf == r_count_24_io_out ? io_r_15_b : _GEN_9794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9796 = 9'h10 == r_count_24_io_out ? io_r_16_b : _GEN_9795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9797 = 9'h11 == r_count_24_io_out ? io_r_17_b : _GEN_9796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9798 = 9'h12 == r_count_24_io_out ? io_r_18_b : _GEN_9797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9799 = 9'h13 == r_count_24_io_out ? io_r_19_b : _GEN_9798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9800 = 9'h14 == r_count_24_io_out ? io_r_20_b : _GEN_9799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9801 = 9'h15 == r_count_24_io_out ? io_r_21_b : _GEN_9800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9802 = 9'h16 == r_count_24_io_out ? io_r_22_b : _GEN_9801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9803 = 9'h17 == r_count_24_io_out ? io_r_23_b : _GEN_9802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9804 = 9'h18 == r_count_24_io_out ? io_r_24_b : _GEN_9803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9805 = 9'h19 == r_count_24_io_out ? io_r_25_b : _GEN_9804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9806 = 9'h1a == r_count_24_io_out ? io_r_26_b : _GEN_9805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9807 = 9'h1b == r_count_24_io_out ? io_r_27_b : _GEN_9806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9808 = 9'h1c == r_count_24_io_out ? io_r_28_b : _GEN_9807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9809 = 9'h1d == r_count_24_io_out ? io_r_29_b : _GEN_9808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9810 = 9'h1e == r_count_24_io_out ? io_r_30_b : _GEN_9809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9811 = 9'h1f == r_count_24_io_out ? io_r_31_b : _GEN_9810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9812 = 9'h20 == r_count_24_io_out ? io_r_32_b : _GEN_9811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9813 = 9'h21 == r_count_24_io_out ? io_r_33_b : _GEN_9812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9814 = 9'h22 == r_count_24_io_out ? io_r_34_b : _GEN_9813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9815 = 9'h23 == r_count_24_io_out ? io_r_35_b : _GEN_9814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9816 = 9'h24 == r_count_24_io_out ? io_r_36_b : _GEN_9815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9817 = 9'h25 == r_count_24_io_out ? io_r_37_b : _GEN_9816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9818 = 9'h26 == r_count_24_io_out ? io_r_38_b : _GEN_9817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9819 = 9'h27 == r_count_24_io_out ? io_r_39_b : _GEN_9818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9820 = 9'h28 == r_count_24_io_out ? io_r_40_b : _GEN_9819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9821 = 9'h29 == r_count_24_io_out ? io_r_41_b : _GEN_9820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9822 = 9'h2a == r_count_24_io_out ? io_r_42_b : _GEN_9821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9823 = 9'h2b == r_count_24_io_out ? io_r_43_b : _GEN_9822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9824 = 9'h2c == r_count_24_io_out ? io_r_44_b : _GEN_9823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9825 = 9'h2d == r_count_24_io_out ? io_r_45_b : _GEN_9824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9826 = 9'h2e == r_count_24_io_out ? io_r_46_b : _GEN_9825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9827 = 9'h2f == r_count_24_io_out ? io_r_47_b : _GEN_9826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9828 = 9'h30 == r_count_24_io_out ? io_r_48_b : _GEN_9827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9829 = 9'h31 == r_count_24_io_out ? io_r_49_b : _GEN_9828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9830 = 9'h32 == r_count_24_io_out ? io_r_50_b : _GEN_9829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9831 = 9'h33 == r_count_24_io_out ? io_r_51_b : _GEN_9830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9832 = 9'h34 == r_count_24_io_out ? io_r_52_b : _GEN_9831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9833 = 9'h35 == r_count_24_io_out ? io_r_53_b : _GEN_9832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9834 = 9'h36 == r_count_24_io_out ? io_r_54_b : _GEN_9833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9835 = 9'h37 == r_count_24_io_out ? io_r_55_b : _GEN_9834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9836 = 9'h38 == r_count_24_io_out ? io_r_56_b : _GEN_9835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9837 = 9'h39 == r_count_24_io_out ? io_r_57_b : _GEN_9836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9838 = 9'h3a == r_count_24_io_out ? io_r_58_b : _GEN_9837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9839 = 9'h3b == r_count_24_io_out ? io_r_59_b : _GEN_9838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9840 = 9'h3c == r_count_24_io_out ? io_r_60_b : _GEN_9839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9841 = 9'h3d == r_count_24_io_out ? io_r_61_b : _GEN_9840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9842 = 9'h3e == r_count_24_io_out ? io_r_62_b : _GEN_9841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9843 = 9'h3f == r_count_24_io_out ? io_r_63_b : _GEN_9842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9844 = 9'h40 == r_count_24_io_out ? io_r_64_b : _GEN_9843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9845 = 9'h41 == r_count_24_io_out ? io_r_65_b : _GEN_9844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9846 = 9'h42 == r_count_24_io_out ? io_r_66_b : _GEN_9845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9847 = 9'h43 == r_count_24_io_out ? io_r_67_b : _GEN_9846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9848 = 9'h44 == r_count_24_io_out ? io_r_68_b : _GEN_9847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9849 = 9'h45 == r_count_24_io_out ? io_r_69_b : _GEN_9848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9850 = 9'h46 == r_count_24_io_out ? io_r_70_b : _GEN_9849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9851 = 9'h47 == r_count_24_io_out ? io_r_71_b : _GEN_9850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9852 = 9'h48 == r_count_24_io_out ? io_r_72_b : _GEN_9851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9853 = 9'h49 == r_count_24_io_out ? io_r_73_b : _GEN_9852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9854 = 9'h4a == r_count_24_io_out ? io_r_74_b : _GEN_9853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9855 = 9'h4b == r_count_24_io_out ? io_r_75_b : _GEN_9854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9856 = 9'h4c == r_count_24_io_out ? io_r_76_b : _GEN_9855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9857 = 9'h4d == r_count_24_io_out ? io_r_77_b : _GEN_9856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9858 = 9'h4e == r_count_24_io_out ? io_r_78_b : _GEN_9857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9859 = 9'h4f == r_count_24_io_out ? io_r_79_b : _GEN_9858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9860 = 9'h50 == r_count_24_io_out ? io_r_80_b : _GEN_9859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9861 = 9'h51 == r_count_24_io_out ? io_r_81_b : _GEN_9860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9862 = 9'h52 == r_count_24_io_out ? io_r_82_b : _GEN_9861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9863 = 9'h53 == r_count_24_io_out ? io_r_83_b : _GEN_9862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9864 = 9'h54 == r_count_24_io_out ? io_r_84_b : _GEN_9863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9865 = 9'h55 == r_count_24_io_out ? io_r_85_b : _GEN_9864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9866 = 9'h56 == r_count_24_io_out ? io_r_86_b : _GEN_9865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9867 = 9'h57 == r_count_24_io_out ? io_r_87_b : _GEN_9866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9868 = 9'h58 == r_count_24_io_out ? io_r_88_b : _GEN_9867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9869 = 9'h59 == r_count_24_io_out ? io_r_89_b : _GEN_9868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9870 = 9'h5a == r_count_24_io_out ? io_r_90_b : _GEN_9869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9871 = 9'h5b == r_count_24_io_out ? io_r_91_b : _GEN_9870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9872 = 9'h5c == r_count_24_io_out ? io_r_92_b : _GEN_9871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9873 = 9'h5d == r_count_24_io_out ? io_r_93_b : _GEN_9872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9874 = 9'h5e == r_count_24_io_out ? io_r_94_b : _GEN_9873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9875 = 9'h5f == r_count_24_io_out ? io_r_95_b : _GEN_9874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9876 = 9'h60 == r_count_24_io_out ? io_r_96_b : _GEN_9875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9877 = 9'h61 == r_count_24_io_out ? io_r_97_b : _GEN_9876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9878 = 9'h62 == r_count_24_io_out ? io_r_98_b : _GEN_9877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9879 = 9'h63 == r_count_24_io_out ? io_r_99_b : _GEN_9878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9880 = 9'h64 == r_count_24_io_out ? io_r_100_b : _GEN_9879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9881 = 9'h65 == r_count_24_io_out ? io_r_101_b : _GEN_9880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9882 = 9'h66 == r_count_24_io_out ? io_r_102_b : _GEN_9881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9883 = 9'h67 == r_count_24_io_out ? io_r_103_b : _GEN_9882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9884 = 9'h68 == r_count_24_io_out ? io_r_104_b : _GEN_9883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9885 = 9'h69 == r_count_24_io_out ? io_r_105_b : _GEN_9884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9886 = 9'h6a == r_count_24_io_out ? io_r_106_b : _GEN_9885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9887 = 9'h6b == r_count_24_io_out ? io_r_107_b : _GEN_9886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9888 = 9'h6c == r_count_24_io_out ? io_r_108_b : _GEN_9887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9889 = 9'h6d == r_count_24_io_out ? io_r_109_b : _GEN_9888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9890 = 9'h6e == r_count_24_io_out ? io_r_110_b : _GEN_9889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9891 = 9'h6f == r_count_24_io_out ? io_r_111_b : _GEN_9890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9892 = 9'h70 == r_count_24_io_out ? io_r_112_b : _GEN_9891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9893 = 9'h71 == r_count_24_io_out ? io_r_113_b : _GEN_9892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9894 = 9'h72 == r_count_24_io_out ? io_r_114_b : _GEN_9893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9895 = 9'h73 == r_count_24_io_out ? io_r_115_b : _GEN_9894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9896 = 9'h74 == r_count_24_io_out ? io_r_116_b : _GEN_9895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9897 = 9'h75 == r_count_24_io_out ? io_r_117_b : _GEN_9896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9898 = 9'h76 == r_count_24_io_out ? io_r_118_b : _GEN_9897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9899 = 9'h77 == r_count_24_io_out ? io_r_119_b : _GEN_9898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9900 = 9'h78 == r_count_24_io_out ? io_r_120_b : _GEN_9899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9901 = 9'h79 == r_count_24_io_out ? io_r_121_b : _GEN_9900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9902 = 9'h7a == r_count_24_io_out ? io_r_122_b : _GEN_9901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9903 = 9'h7b == r_count_24_io_out ? io_r_123_b : _GEN_9902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9904 = 9'h7c == r_count_24_io_out ? io_r_124_b : _GEN_9903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9905 = 9'h7d == r_count_24_io_out ? io_r_125_b : _GEN_9904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9906 = 9'h7e == r_count_24_io_out ? io_r_126_b : _GEN_9905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9907 = 9'h7f == r_count_24_io_out ? io_r_127_b : _GEN_9906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9908 = 9'h80 == r_count_24_io_out ? io_r_128_b : _GEN_9907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9909 = 9'h81 == r_count_24_io_out ? io_r_129_b : _GEN_9908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9910 = 9'h82 == r_count_24_io_out ? io_r_130_b : _GEN_9909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9911 = 9'h83 == r_count_24_io_out ? io_r_131_b : _GEN_9910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9912 = 9'h84 == r_count_24_io_out ? io_r_132_b : _GEN_9911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9913 = 9'h85 == r_count_24_io_out ? io_r_133_b : _GEN_9912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9914 = 9'h86 == r_count_24_io_out ? io_r_134_b : _GEN_9913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9915 = 9'h87 == r_count_24_io_out ? io_r_135_b : _GEN_9914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9916 = 9'h88 == r_count_24_io_out ? io_r_136_b : _GEN_9915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9917 = 9'h89 == r_count_24_io_out ? io_r_137_b : _GEN_9916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9918 = 9'h8a == r_count_24_io_out ? io_r_138_b : _GEN_9917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9919 = 9'h8b == r_count_24_io_out ? io_r_139_b : _GEN_9918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9920 = 9'h8c == r_count_24_io_out ? io_r_140_b : _GEN_9919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9921 = 9'h8d == r_count_24_io_out ? io_r_141_b : _GEN_9920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9922 = 9'h8e == r_count_24_io_out ? io_r_142_b : _GEN_9921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9923 = 9'h8f == r_count_24_io_out ? io_r_143_b : _GEN_9922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9924 = 9'h90 == r_count_24_io_out ? io_r_144_b : _GEN_9923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9925 = 9'h91 == r_count_24_io_out ? io_r_145_b : _GEN_9924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9926 = 9'h92 == r_count_24_io_out ? io_r_146_b : _GEN_9925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9927 = 9'h93 == r_count_24_io_out ? io_r_147_b : _GEN_9926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9928 = 9'h94 == r_count_24_io_out ? io_r_148_b : _GEN_9927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9929 = 9'h95 == r_count_24_io_out ? io_r_149_b : _GEN_9928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9930 = 9'h96 == r_count_24_io_out ? io_r_150_b : _GEN_9929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9931 = 9'h97 == r_count_24_io_out ? io_r_151_b : _GEN_9930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9932 = 9'h98 == r_count_24_io_out ? io_r_152_b : _GEN_9931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9933 = 9'h99 == r_count_24_io_out ? io_r_153_b : _GEN_9932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9934 = 9'h9a == r_count_24_io_out ? io_r_154_b : _GEN_9933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9935 = 9'h9b == r_count_24_io_out ? io_r_155_b : _GEN_9934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9936 = 9'h9c == r_count_24_io_out ? io_r_156_b : _GEN_9935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9937 = 9'h9d == r_count_24_io_out ? io_r_157_b : _GEN_9936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9938 = 9'h9e == r_count_24_io_out ? io_r_158_b : _GEN_9937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9939 = 9'h9f == r_count_24_io_out ? io_r_159_b : _GEN_9938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9940 = 9'ha0 == r_count_24_io_out ? io_r_160_b : _GEN_9939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9941 = 9'ha1 == r_count_24_io_out ? io_r_161_b : _GEN_9940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9942 = 9'ha2 == r_count_24_io_out ? io_r_162_b : _GEN_9941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9943 = 9'ha3 == r_count_24_io_out ? io_r_163_b : _GEN_9942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9944 = 9'ha4 == r_count_24_io_out ? io_r_164_b : _GEN_9943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9945 = 9'ha5 == r_count_24_io_out ? io_r_165_b : _GEN_9944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9946 = 9'ha6 == r_count_24_io_out ? io_r_166_b : _GEN_9945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9947 = 9'ha7 == r_count_24_io_out ? io_r_167_b : _GEN_9946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9948 = 9'ha8 == r_count_24_io_out ? io_r_168_b : _GEN_9947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9949 = 9'ha9 == r_count_24_io_out ? io_r_169_b : _GEN_9948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9950 = 9'haa == r_count_24_io_out ? io_r_170_b : _GEN_9949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9951 = 9'hab == r_count_24_io_out ? io_r_171_b : _GEN_9950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9952 = 9'hac == r_count_24_io_out ? io_r_172_b : _GEN_9951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9953 = 9'had == r_count_24_io_out ? io_r_173_b : _GEN_9952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9954 = 9'hae == r_count_24_io_out ? io_r_174_b : _GEN_9953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9955 = 9'haf == r_count_24_io_out ? io_r_175_b : _GEN_9954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9956 = 9'hb0 == r_count_24_io_out ? io_r_176_b : _GEN_9955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9957 = 9'hb1 == r_count_24_io_out ? io_r_177_b : _GEN_9956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9958 = 9'hb2 == r_count_24_io_out ? io_r_178_b : _GEN_9957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9959 = 9'hb3 == r_count_24_io_out ? io_r_179_b : _GEN_9958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9960 = 9'hb4 == r_count_24_io_out ? io_r_180_b : _GEN_9959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9961 = 9'hb5 == r_count_24_io_out ? io_r_181_b : _GEN_9960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9962 = 9'hb6 == r_count_24_io_out ? io_r_182_b : _GEN_9961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9963 = 9'hb7 == r_count_24_io_out ? io_r_183_b : _GEN_9962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9964 = 9'hb8 == r_count_24_io_out ? io_r_184_b : _GEN_9963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9965 = 9'hb9 == r_count_24_io_out ? io_r_185_b : _GEN_9964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9966 = 9'hba == r_count_24_io_out ? io_r_186_b : _GEN_9965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9967 = 9'hbb == r_count_24_io_out ? io_r_187_b : _GEN_9966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9968 = 9'hbc == r_count_24_io_out ? io_r_188_b : _GEN_9967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9969 = 9'hbd == r_count_24_io_out ? io_r_189_b : _GEN_9968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9970 = 9'hbe == r_count_24_io_out ? io_r_190_b : _GEN_9969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9971 = 9'hbf == r_count_24_io_out ? io_r_191_b : _GEN_9970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9972 = 9'hc0 == r_count_24_io_out ? io_r_192_b : _GEN_9971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9973 = 9'hc1 == r_count_24_io_out ? io_r_193_b : _GEN_9972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9974 = 9'hc2 == r_count_24_io_out ? io_r_194_b : _GEN_9973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9975 = 9'hc3 == r_count_24_io_out ? io_r_195_b : _GEN_9974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9976 = 9'hc4 == r_count_24_io_out ? io_r_196_b : _GEN_9975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9977 = 9'hc5 == r_count_24_io_out ? io_r_197_b : _GEN_9976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9978 = 9'hc6 == r_count_24_io_out ? io_r_198_b : _GEN_9977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9979 = 9'hc7 == r_count_24_io_out ? io_r_199_b : _GEN_9978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9980 = 9'hc8 == r_count_24_io_out ? io_r_200_b : _GEN_9979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9981 = 9'hc9 == r_count_24_io_out ? io_r_201_b : _GEN_9980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9982 = 9'hca == r_count_24_io_out ? io_r_202_b : _GEN_9981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9983 = 9'hcb == r_count_24_io_out ? io_r_203_b : _GEN_9982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9984 = 9'hcc == r_count_24_io_out ? io_r_204_b : _GEN_9983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9985 = 9'hcd == r_count_24_io_out ? io_r_205_b : _GEN_9984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9986 = 9'hce == r_count_24_io_out ? io_r_206_b : _GEN_9985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9987 = 9'hcf == r_count_24_io_out ? io_r_207_b : _GEN_9986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9988 = 9'hd0 == r_count_24_io_out ? io_r_208_b : _GEN_9987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9989 = 9'hd1 == r_count_24_io_out ? io_r_209_b : _GEN_9988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9990 = 9'hd2 == r_count_24_io_out ? io_r_210_b : _GEN_9989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9991 = 9'hd3 == r_count_24_io_out ? io_r_211_b : _GEN_9990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9992 = 9'hd4 == r_count_24_io_out ? io_r_212_b : _GEN_9991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9993 = 9'hd5 == r_count_24_io_out ? io_r_213_b : _GEN_9992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9994 = 9'hd6 == r_count_24_io_out ? io_r_214_b : _GEN_9993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9995 = 9'hd7 == r_count_24_io_out ? io_r_215_b : _GEN_9994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9996 = 9'hd8 == r_count_24_io_out ? io_r_216_b : _GEN_9995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9997 = 9'hd9 == r_count_24_io_out ? io_r_217_b : _GEN_9996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9998 = 9'hda == r_count_24_io_out ? io_r_218_b : _GEN_9997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9999 = 9'hdb == r_count_24_io_out ? io_r_219_b : _GEN_9998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10000 = 9'hdc == r_count_24_io_out ? io_r_220_b : _GEN_9999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10001 = 9'hdd == r_count_24_io_out ? io_r_221_b : _GEN_10000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10002 = 9'hde == r_count_24_io_out ? io_r_222_b : _GEN_10001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10003 = 9'hdf == r_count_24_io_out ? io_r_223_b : _GEN_10002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10004 = 9'he0 == r_count_24_io_out ? io_r_224_b : _GEN_10003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10005 = 9'he1 == r_count_24_io_out ? io_r_225_b : _GEN_10004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10006 = 9'he2 == r_count_24_io_out ? io_r_226_b : _GEN_10005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10007 = 9'he3 == r_count_24_io_out ? io_r_227_b : _GEN_10006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10008 = 9'he4 == r_count_24_io_out ? io_r_228_b : _GEN_10007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10009 = 9'he5 == r_count_24_io_out ? io_r_229_b : _GEN_10008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10010 = 9'he6 == r_count_24_io_out ? io_r_230_b : _GEN_10009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10011 = 9'he7 == r_count_24_io_out ? io_r_231_b : _GEN_10010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10012 = 9'he8 == r_count_24_io_out ? io_r_232_b : _GEN_10011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10013 = 9'he9 == r_count_24_io_out ? io_r_233_b : _GEN_10012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10014 = 9'hea == r_count_24_io_out ? io_r_234_b : _GEN_10013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10015 = 9'heb == r_count_24_io_out ? io_r_235_b : _GEN_10014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10016 = 9'hec == r_count_24_io_out ? io_r_236_b : _GEN_10015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10017 = 9'hed == r_count_24_io_out ? io_r_237_b : _GEN_10016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10018 = 9'hee == r_count_24_io_out ? io_r_238_b : _GEN_10017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10019 = 9'hef == r_count_24_io_out ? io_r_239_b : _GEN_10018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10020 = 9'hf0 == r_count_24_io_out ? io_r_240_b : _GEN_10019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10021 = 9'hf1 == r_count_24_io_out ? io_r_241_b : _GEN_10020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10022 = 9'hf2 == r_count_24_io_out ? io_r_242_b : _GEN_10021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10023 = 9'hf3 == r_count_24_io_out ? io_r_243_b : _GEN_10022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10024 = 9'hf4 == r_count_24_io_out ? io_r_244_b : _GEN_10023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10025 = 9'hf5 == r_count_24_io_out ? io_r_245_b : _GEN_10024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10026 = 9'hf6 == r_count_24_io_out ? io_r_246_b : _GEN_10025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10027 = 9'hf7 == r_count_24_io_out ? io_r_247_b : _GEN_10026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10028 = 9'hf8 == r_count_24_io_out ? io_r_248_b : _GEN_10027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10029 = 9'hf9 == r_count_24_io_out ? io_r_249_b : _GEN_10028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10030 = 9'hfa == r_count_24_io_out ? io_r_250_b : _GEN_10029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10031 = 9'hfb == r_count_24_io_out ? io_r_251_b : _GEN_10030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10032 = 9'hfc == r_count_24_io_out ? io_r_252_b : _GEN_10031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10033 = 9'hfd == r_count_24_io_out ? io_r_253_b : _GEN_10032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10034 = 9'hfe == r_count_24_io_out ? io_r_254_b : _GEN_10033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10035 = 9'hff == r_count_24_io_out ? io_r_255_b : _GEN_10034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10036 = 9'h100 == r_count_24_io_out ? io_r_256_b : _GEN_10035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10037 = 9'h101 == r_count_24_io_out ? io_r_257_b : _GEN_10036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10038 = 9'h102 == r_count_24_io_out ? io_r_258_b : _GEN_10037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10039 = 9'h103 == r_count_24_io_out ? io_r_259_b : _GEN_10038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10040 = 9'h104 == r_count_24_io_out ? io_r_260_b : _GEN_10039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10041 = 9'h105 == r_count_24_io_out ? io_r_261_b : _GEN_10040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10042 = 9'h106 == r_count_24_io_out ? io_r_262_b : _GEN_10041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10043 = 9'h107 == r_count_24_io_out ? io_r_263_b : _GEN_10042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10044 = 9'h108 == r_count_24_io_out ? io_r_264_b : _GEN_10043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10045 = 9'h109 == r_count_24_io_out ? io_r_265_b : _GEN_10044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10046 = 9'h10a == r_count_24_io_out ? io_r_266_b : _GEN_10045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10047 = 9'h10b == r_count_24_io_out ? io_r_267_b : _GEN_10046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10048 = 9'h10c == r_count_24_io_out ? io_r_268_b : _GEN_10047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10049 = 9'h10d == r_count_24_io_out ? io_r_269_b : _GEN_10048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10050 = 9'h10e == r_count_24_io_out ? io_r_270_b : _GEN_10049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10051 = 9'h10f == r_count_24_io_out ? io_r_271_b : _GEN_10050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10052 = 9'h110 == r_count_24_io_out ? io_r_272_b : _GEN_10051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10053 = 9'h111 == r_count_24_io_out ? io_r_273_b : _GEN_10052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10054 = 9'h112 == r_count_24_io_out ? io_r_274_b : _GEN_10053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10055 = 9'h113 == r_count_24_io_out ? io_r_275_b : _GEN_10054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10056 = 9'h114 == r_count_24_io_out ? io_r_276_b : _GEN_10055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10057 = 9'h115 == r_count_24_io_out ? io_r_277_b : _GEN_10056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10058 = 9'h116 == r_count_24_io_out ? io_r_278_b : _GEN_10057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10059 = 9'h117 == r_count_24_io_out ? io_r_279_b : _GEN_10058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10060 = 9'h118 == r_count_24_io_out ? io_r_280_b : _GEN_10059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10061 = 9'h119 == r_count_24_io_out ? io_r_281_b : _GEN_10060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10062 = 9'h11a == r_count_24_io_out ? io_r_282_b : _GEN_10061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10063 = 9'h11b == r_count_24_io_out ? io_r_283_b : _GEN_10062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10064 = 9'h11c == r_count_24_io_out ? io_r_284_b : _GEN_10063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10065 = 9'h11d == r_count_24_io_out ? io_r_285_b : _GEN_10064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10066 = 9'h11e == r_count_24_io_out ? io_r_286_b : _GEN_10065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10067 = 9'h11f == r_count_24_io_out ? io_r_287_b : _GEN_10066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10068 = 9'h120 == r_count_24_io_out ? io_r_288_b : _GEN_10067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10069 = 9'h121 == r_count_24_io_out ? io_r_289_b : _GEN_10068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10070 = 9'h122 == r_count_24_io_out ? io_r_290_b : _GEN_10069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10071 = 9'h123 == r_count_24_io_out ? io_r_291_b : _GEN_10070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10072 = 9'h124 == r_count_24_io_out ? io_r_292_b : _GEN_10071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10073 = 9'h125 == r_count_24_io_out ? io_r_293_b : _GEN_10072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10074 = 9'h126 == r_count_24_io_out ? io_r_294_b : _GEN_10073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10075 = 9'h127 == r_count_24_io_out ? io_r_295_b : _GEN_10074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10076 = 9'h128 == r_count_24_io_out ? io_r_296_b : _GEN_10075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10077 = 9'h129 == r_count_24_io_out ? io_r_297_b : _GEN_10076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10078 = 9'h12a == r_count_24_io_out ? io_r_298_b : _GEN_10077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10079 = 9'h12b == r_count_24_io_out ? io_r_299_b : _GEN_10078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10080 = 9'h12c == r_count_24_io_out ? io_r_300_b : _GEN_10079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10081 = 9'h12d == r_count_24_io_out ? io_r_301_b : _GEN_10080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10082 = 9'h12e == r_count_24_io_out ? io_r_302_b : _GEN_10081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10083 = 9'h12f == r_count_24_io_out ? io_r_303_b : _GEN_10082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10084 = 9'h130 == r_count_24_io_out ? io_r_304_b : _GEN_10083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10085 = 9'h131 == r_count_24_io_out ? io_r_305_b : _GEN_10084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10086 = 9'h132 == r_count_24_io_out ? io_r_306_b : _GEN_10085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10087 = 9'h133 == r_count_24_io_out ? io_r_307_b : _GEN_10086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10088 = 9'h134 == r_count_24_io_out ? io_r_308_b : _GEN_10087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10089 = 9'h135 == r_count_24_io_out ? io_r_309_b : _GEN_10088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10090 = 9'h136 == r_count_24_io_out ? io_r_310_b : _GEN_10089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10091 = 9'h137 == r_count_24_io_out ? io_r_311_b : _GEN_10090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10092 = 9'h138 == r_count_24_io_out ? io_r_312_b : _GEN_10091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10093 = 9'h139 == r_count_24_io_out ? io_r_313_b : _GEN_10092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10094 = 9'h13a == r_count_24_io_out ? io_r_314_b : _GEN_10093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10095 = 9'h13b == r_count_24_io_out ? io_r_315_b : _GEN_10094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10096 = 9'h13c == r_count_24_io_out ? io_r_316_b : _GEN_10095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10097 = 9'h13d == r_count_24_io_out ? io_r_317_b : _GEN_10096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10098 = 9'h13e == r_count_24_io_out ? io_r_318_b : _GEN_10097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10099 = 9'h13f == r_count_24_io_out ? io_r_319_b : _GEN_10098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10100 = 9'h140 == r_count_24_io_out ? io_r_320_b : _GEN_10099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10101 = 9'h141 == r_count_24_io_out ? io_r_321_b : _GEN_10100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10102 = 9'h142 == r_count_24_io_out ? io_r_322_b : _GEN_10101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10103 = 9'h143 == r_count_24_io_out ? io_r_323_b : _GEN_10102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10104 = 9'h144 == r_count_24_io_out ? io_r_324_b : _GEN_10103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10105 = 9'h145 == r_count_24_io_out ? io_r_325_b : _GEN_10104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10106 = 9'h146 == r_count_24_io_out ? io_r_326_b : _GEN_10105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10107 = 9'h147 == r_count_24_io_out ? io_r_327_b : _GEN_10106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10108 = 9'h148 == r_count_24_io_out ? io_r_328_b : _GEN_10107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10109 = 9'h149 == r_count_24_io_out ? io_r_329_b : _GEN_10108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10110 = 9'h14a == r_count_24_io_out ? io_r_330_b : _GEN_10109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10111 = 9'h14b == r_count_24_io_out ? io_r_331_b : _GEN_10110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10112 = 9'h14c == r_count_24_io_out ? io_r_332_b : _GEN_10111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10113 = 9'h14d == r_count_24_io_out ? io_r_333_b : _GEN_10112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10114 = 9'h14e == r_count_24_io_out ? io_r_334_b : _GEN_10113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10115 = 9'h14f == r_count_24_io_out ? io_r_335_b : _GEN_10114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10116 = 9'h150 == r_count_24_io_out ? io_r_336_b : _GEN_10115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10117 = 9'h151 == r_count_24_io_out ? io_r_337_b : _GEN_10116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10118 = 9'h152 == r_count_24_io_out ? io_r_338_b : _GEN_10117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10119 = 9'h153 == r_count_24_io_out ? io_r_339_b : _GEN_10118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10120 = 9'h154 == r_count_24_io_out ? io_r_340_b : _GEN_10119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10121 = 9'h155 == r_count_24_io_out ? io_r_341_b : _GEN_10120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10122 = 9'h156 == r_count_24_io_out ? io_r_342_b : _GEN_10121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10123 = 9'h157 == r_count_24_io_out ? io_r_343_b : _GEN_10122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10124 = 9'h158 == r_count_24_io_out ? io_r_344_b : _GEN_10123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10125 = 9'h159 == r_count_24_io_out ? io_r_345_b : _GEN_10124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10126 = 9'h15a == r_count_24_io_out ? io_r_346_b : _GEN_10125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10127 = 9'h15b == r_count_24_io_out ? io_r_347_b : _GEN_10126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10128 = 9'h15c == r_count_24_io_out ? io_r_348_b : _GEN_10127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10129 = 9'h15d == r_count_24_io_out ? io_r_349_b : _GEN_10128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10130 = 9'h15e == r_count_24_io_out ? io_r_350_b : _GEN_10129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10131 = 9'h15f == r_count_24_io_out ? io_r_351_b : _GEN_10130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10132 = 9'h160 == r_count_24_io_out ? io_r_352_b : _GEN_10131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10133 = 9'h161 == r_count_24_io_out ? io_r_353_b : _GEN_10132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10134 = 9'h162 == r_count_24_io_out ? io_r_354_b : _GEN_10133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10135 = 9'h163 == r_count_24_io_out ? io_r_355_b : _GEN_10134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10136 = 9'h164 == r_count_24_io_out ? io_r_356_b : _GEN_10135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10137 = 9'h165 == r_count_24_io_out ? io_r_357_b : _GEN_10136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10138 = 9'h166 == r_count_24_io_out ? io_r_358_b : _GEN_10137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10139 = 9'h167 == r_count_24_io_out ? io_r_359_b : _GEN_10138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10140 = 9'h168 == r_count_24_io_out ? io_r_360_b : _GEN_10139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10141 = 9'h169 == r_count_24_io_out ? io_r_361_b : _GEN_10140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10142 = 9'h16a == r_count_24_io_out ? io_r_362_b : _GEN_10141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10143 = 9'h16b == r_count_24_io_out ? io_r_363_b : _GEN_10142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10144 = 9'h16c == r_count_24_io_out ? io_r_364_b : _GEN_10143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10145 = 9'h16d == r_count_24_io_out ? io_r_365_b : _GEN_10144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10146 = 9'h16e == r_count_24_io_out ? io_r_366_b : _GEN_10145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10147 = 9'h16f == r_count_24_io_out ? io_r_367_b : _GEN_10146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10148 = 9'h170 == r_count_24_io_out ? io_r_368_b : _GEN_10147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10149 = 9'h171 == r_count_24_io_out ? io_r_369_b : _GEN_10148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10150 = 9'h172 == r_count_24_io_out ? io_r_370_b : _GEN_10149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10151 = 9'h173 == r_count_24_io_out ? io_r_371_b : _GEN_10150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10152 = 9'h174 == r_count_24_io_out ? io_r_372_b : _GEN_10151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10153 = 9'h175 == r_count_24_io_out ? io_r_373_b : _GEN_10152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10154 = 9'h176 == r_count_24_io_out ? io_r_374_b : _GEN_10153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10155 = 9'h177 == r_count_24_io_out ? io_r_375_b : _GEN_10154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10156 = 9'h178 == r_count_24_io_out ? io_r_376_b : _GEN_10155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10157 = 9'h179 == r_count_24_io_out ? io_r_377_b : _GEN_10156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10158 = 9'h17a == r_count_24_io_out ? io_r_378_b : _GEN_10157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10159 = 9'h17b == r_count_24_io_out ? io_r_379_b : _GEN_10158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10160 = 9'h17c == r_count_24_io_out ? io_r_380_b : _GEN_10159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10161 = 9'h17d == r_count_24_io_out ? io_r_381_b : _GEN_10160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10162 = 9'h17e == r_count_24_io_out ? io_r_382_b : _GEN_10161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10163 = 9'h17f == r_count_24_io_out ? io_r_383_b : _GEN_10162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10164 = 9'h180 == r_count_24_io_out ? io_r_384_b : _GEN_10163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10165 = 9'h181 == r_count_24_io_out ? io_r_385_b : _GEN_10164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10166 = 9'h182 == r_count_24_io_out ? io_r_386_b : _GEN_10165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10167 = 9'h183 == r_count_24_io_out ? io_r_387_b : _GEN_10166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10168 = 9'h184 == r_count_24_io_out ? io_r_388_b : _GEN_10167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10169 = 9'h185 == r_count_24_io_out ? io_r_389_b : _GEN_10168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10170 = 9'h186 == r_count_24_io_out ? io_r_390_b : _GEN_10169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10171 = 9'h187 == r_count_24_io_out ? io_r_391_b : _GEN_10170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10172 = 9'h188 == r_count_24_io_out ? io_r_392_b : _GEN_10171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10173 = 9'h189 == r_count_24_io_out ? io_r_393_b : _GEN_10172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10174 = 9'h18a == r_count_24_io_out ? io_r_394_b : _GEN_10173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10175 = 9'h18b == r_count_24_io_out ? io_r_395_b : _GEN_10174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10176 = 9'h18c == r_count_24_io_out ? io_r_396_b : _GEN_10175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10177 = 9'h18d == r_count_24_io_out ? io_r_397_b : _GEN_10176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10178 = 9'h18e == r_count_24_io_out ? io_r_398_b : _GEN_10177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10181 = 9'h1 == r_count_25_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10182 = 9'h2 == r_count_25_io_out ? io_r_2_b : _GEN_10181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10183 = 9'h3 == r_count_25_io_out ? io_r_3_b : _GEN_10182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10184 = 9'h4 == r_count_25_io_out ? io_r_4_b : _GEN_10183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10185 = 9'h5 == r_count_25_io_out ? io_r_5_b : _GEN_10184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10186 = 9'h6 == r_count_25_io_out ? io_r_6_b : _GEN_10185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10187 = 9'h7 == r_count_25_io_out ? io_r_7_b : _GEN_10186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10188 = 9'h8 == r_count_25_io_out ? io_r_8_b : _GEN_10187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10189 = 9'h9 == r_count_25_io_out ? io_r_9_b : _GEN_10188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10190 = 9'ha == r_count_25_io_out ? io_r_10_b : _GEN_10189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10191 = 9'hb == r_count_25_io_out ? io_r_11_b : _GEN_10190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10192 = 9'hc == r_count_25_io_out ? io_r_12_b : _GEN_10191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10193 = 9'hd == r_count_25_io_out ? io_r_13_b : _GEN_10192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10194 = 9'he == r_count_25_io_out ? io_r_14_b : _GEN_10193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10195 = 9'hf == r_count_25_io_out ? io_r_15_b : _GEN_10194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10196 = 9'h10 == r_count_25_io_out ? io_r_16_b : _GEN_10195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10197 = 9'h11 == r_count_25_io_out ? io_r_17_b : _GEN_10196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10198 = 9'h12 == r_count_25_io_out ? io_r_18_b : _GEN_10197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10199 = 9'h13 == r_count_25_io_out ? io_r_19_b : _GEN_10198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10200 = 9'h14 == r_count_25_io_out ? io_r_20_b : _GEN_10199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10201 = 9'h15 == r_count_25_io_out ? io_r_21_b : _GEN_10200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10202 = 9'h16 == r_count_25_io_out ? io_r_22_b : _GEN_10201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10203 = 9'h17 == r_count_25_io_out ? io_r_23_b : _GEN_10202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10204 = 9'h18 == r_count_25_io_out ? io_r_24_b : _GEN_10203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10205 = 9'h19 == r_count_25_io_out ? io_r_25_b : _GEN_10204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10206 = 9'h1a == r_count_25_io_out ? io_r_26_b : _GEN_10205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10207 = 9'h1b == r_count_25_io_out ? io_r_27_b : _GEN_10206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10208 = 9'h1c == r_count_25_io_out ? io_r_28_b : _GEN_10207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10209 = 9'h1d == r_count_25_io_out ? io_r_29_b : _GEN_10208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10210 = 9'h1e == r_count_25_io_out ? io_r_30_b : _GEN_10209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10211 = 9'h1f == r_count_25_io_out ? io_r_31_b : _GEN_10210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10212 = 9'h20 == r_count_25_io_out ? io_r_32_b : _GEN_10211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10213 = 9'h21 == r_count_25_io_out ? io_r_33_b : _GEN_10212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10214 = 9'h22 == r_count_25_io_out ? io_r_34_b : _GEN_10213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10215 = 9'h23 == r_count_25_io_out ? io_r_35_b : _GEN_10214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10216 = 9'h24 == r_count_25_io_out ? io_r_36_b : _GEN_10215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10217 = 9'h25 == r_count_25_io_out ? io_r_37_b : _GEN_10216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10218 = 9'h26 == r_count_25_io_out ? io_r_38_b : _GEN_10217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10219 = 9'h27 == r_count_25_io_out ? io_r_39_b : _GEN_10218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10220 = 9'h28 == r_count_25_io_out ? io_r_40_b : _GEN_10219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10221 = 9'h29 == r_count_25_io_out ? io_r_41_b : _GEN_10220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10222 = 9'h2a == r_count_25_io_out ? io_r_42_b : _GEN_10221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10223 = 9'h2b == r_count_25_io_out ? io_r_43_b : _GEN_10222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10224 = 9'h2c == r_count_25_io_out ? io_r_44_b : _GEN_10223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10225 = 9'h2d == r_count_25_io_out ? io_r_45_b : _GEN_10224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10226 = 9'h2e == r_count_25_io_out ? io_r_46_b : _GEN_10225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10227 = 9'h2f == r_count_25_io_out ? io_r_47_b : _GEN_10226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10228 = 9'h30 == r_count_25_io_out ? io_r_48_b : _GEN_10227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10229 = 9'h31 == r_count_25_io_out ? io_r_49_b : _GEN_10228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10230 = 9'h32 == r_count_25_io_out ? io_r_50_b : _GEN_10229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10231 = 9'h33 == r_count_25_io_out ? io_r_51_b : _GEN_10230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10232 = 9'h34 == r_count_25_io_out ? io_r_52_b : _GEN_10231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10233 = 9'h35 == r_count_25_io_out ? io_r_53_b : _GEN_10232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10234 = 9'h36 == r_count_25_io_out ? io_r_54_b : _GEN_10233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10235 = 9'h37 == r_count_25_io_out ? io_r_55_b : _GEN_10234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10236 = 9'h38 == r_count_25_io_out ? io_r_56_b : _GEN_10235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10237 = 9'h39 == r_count_25_io_out ? io_r_57_b : _GEN_10236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10238 = 9'h3a == r_count_25_io_out ? io_r_58_b : _GEN_10237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10239 = 9'h3b == r_count_25_io_out ? io_r_59_b : _GEN_10238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10240 = 9'h3c == r_count_25_io_out ? io_r_60_b : _GEN_10239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10241 = 9'h3d == r_count_25_io_out ? io_r_61_b : _GEN_10240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10242 = 9'h3e == r_count_25_io_out ? io_r_62_b : _GEN_10241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10243 = 9'h3f == r_count_25_io_out ? io_r_63_b : _GEN_10242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10244 = 9'h40 == r_count_25_io_out ? io_r_64_b : _GEN_10243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10245 = 9'h41 == r_count_25_io_out ? io_r_65_b : _GEN_10244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10246 = 9'h42 == r_count_25_io_out ? io_r_66_b : _GEN_10245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10247 = 9'h43 == r_count_25_io_out ? io_r_67_b : _GEN_10246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10248 = 9'h44 == r_count_25_io_out ? io_r_68_b : _GEN_10247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10249 = 9'h45 == r_count_25_io_out ? io_r_69_b : _GEN_10248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10250 = 9'h46 == r_count_25_io_out ? io_r_70_b : _GEN_10249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10251 = 9'h47 == r_count_25_io_out ? io_r_71_b : _GEN_10250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10252 = 9'h48 == r_count_25_io_out ? io_r_72_b : _GEN_10251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10253 = 9'h49 == r_count_25_io_out ? io_r_73_b : _GEN_10252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10254 = 9'h4a == r_count_25_io_out ? io_r_74_b : _GEN_10253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10255 = 9'h4b == r_count_25_io_out ? io_r_75_b : _GEN_10254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10256 = 9'h4c == r_count_25_io_out ? io_r_76_b : _GEN_10255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10257 = 9'h4d == r_count_25_io_out ? io_r_77_b : _GEN_10256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10258 = 9'h4e == r_count_25_io_out ? io_r_78_b : _GEN_10257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10259 = 9'h4f == r_count_25_io_out ? io_r_79_b : _GEN_10258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10260 = 9'h50 == r_count_25_io_out ? io_r_80_b : _GEN_10259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10261 = 9'h51 == r_count_25_io_out ? io_r_81_b : _GEN_10260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10262 = 9'h52 == r_count_25_io_out ? io_r_82_b : _GEN_10261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10263 = 9'h53 == r_count_25_io_out ? io_r_83_b : _GEN_10262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10264 = 9'h54 == r_count_25_io_out ? io_r_84_b : _GEN_10263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10265 = 9'h55 == r_count_25_io_out ? io_r_85_b : _GEN_10264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10266 = 9'h56 == r_count_25_io_out ? io_r_86_b : _GEN_10265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10267 = 9'h57 == r_count_25_io_out ? io_r_87_b : _GEN_10266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10268 = 9'h58 == r_count_25_io_out ? io_r_88_b : _GEN_10267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10269 = 9'h59 == r_count_25_io_out ? io_r_89_b : _GEN_10268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10270 = 9'h5a == r_count_25_io_out ? io_r_90_b : _GEN_10269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10271 = 9'h5b == r_count_25_io_out ? io_r_91_b : _GEN_10270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10272 = 9'h5c == r_count_25_io_out ? io_r_92_b : _GEN_10271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10273 = 9'h5d == r_count_25_io_out ? io_r_93_b : _GEN_10272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10274 = 9'h5e == r_count_25_io_out ? io_r_94_b : _GEN_10273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10275 = 9'h5f == r_count_25_io_out ? io_r_95_b : _GEN_10274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10276 = 9'h60 == r_count_25_io_out ? io_r_96_b : _GEN_10275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10277 = 9'h61 == r_count_25_io_out ? io_r_97_b : _GEN_10276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10278 = 9'h62 == r_count_25_io_out ? io_r_98_b : _GEN_10277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10279 = 9'h63 == r_count_25_io_out ? io_r_99_b : _GEN_10278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10280 = 9'h64 == r_count_25_io_out ? io_r_100_b : _GEN_10279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10281 = 9'h65 == r_count_25_io_out ? io_r_101_b : _GEN_10280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10282 = 9'h66 == r_count_25_io_out ? io_r_102_b : _GEN_10281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10283 = 9'h67 == r_count_25_io_out ? io_r_103_b : _GEN_10282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10284 = 9'h68 == r_count_25_io_out ? io_r_104_b : _GEN_10283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10285 = 9'h69 == r_count_25_io_out ? io_r_105_b : _GEN_10284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10286 = 9'h6a == r_count_25_io_out ? io_r_106_b : _GEN_10285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10287 = 9'h6b == r_count_25_io_out ? io_r_107_b : _GEN_10286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10288 = 9'h6c == r_count_25_io_out ? io_r_108_b : _GEN_10287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10289 = 9'h6d == r_count_25_io_out ? io_r_109_b : _GEN_10288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10290 = 9'h6e == r_count_25_io_out ? io_r_110_b : _GEN_10289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10291 = 9'h6f == r_count_25_io_out ? io_r_111_b : _GEN_10290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10292 = 9'h70 == r_count_25_io_out ? io_r_112_b : _GEN_10291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10293 = 9'h71 == r_count_25_io_out ? io_r_113_b : _GEN_10292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10294 = 9'h72 == r_count_25_io_out ? io_r_114_b : _GEN_10293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10295 = 9'h73 == r_count_25_io_out ? io_r_115_b : _GEN_10294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10296 = 9'h74 == r_count_25_io_out ? io_r_116_b : _GEN_10295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10297 = 9'h75 == r_count_25_io_out ? io_r_117_b : _GEN_10296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10298 = 9'h76 == r_count_25_io_out ? io_r_118_b : _GEN_10297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10299 = 9'h77 == r_count_25_io_out ? io_r_119_b : _GEN_10298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10300 = 9'h78 == r_count_25_io_out ? io_r_120_b : _GEN_10299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10301 = 9'h79 == r_count_25_io_out ? io_r_121_b : _GEN_10300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10302 = 9'h7a == r_count_25_io_out ? io_r_122_b : _GEN_10301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10303 = 9'h7b == r_count_25_io_out ? io_r_123_b : _GEN_10302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10304 = 9'h7c == r_count_25_io_out ? io_r_124_b : _GEN_10303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10305 = 9'h7d == r_count_25_io_out ? io_r_125_b : _GEN_10304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10306 = 9'h7e == r_count_25_io_out ? io_r_126_b : _GEN_10305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10307 = 9'h7f == r_count_25_io_out ? io_r_127_b : _GEN_10306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10308 = 9'h80 == r_count_25_io_out ? io_r_128_b : _GEN_10307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10309 = 9'h81 == r_count_25_io_out ? io_r_129_b : _GEN_10308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10310 = 9'h82 == r_count_25_io_out ? io_r_130_b : _GEN_10309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10311 = 9'h83 == r_count_25_io_out ? io_r_131_b : _GEN_10310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10312 = 9'h84 == r_count_25_io_out ? io_r_132_b : _GEN_10311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10313 = 9'h85 == r_count_25_io_out ? io_r_133_b : _GEN_10312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10314 = 9'h86 == r_count_25_io_out ? io_r_134_b : _GEN_10313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10315 = 9'h87 == r_count_25_io_out ? io_r_135_b : _GEN_10314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10316 = 9'h88 == r_count_25_io_out ? io_r_136_b : _GEN_10315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10317 = 9'h89 == r_count_25_io_out ? io_r_137_b : _GEN_10316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10318 = 9'h8a == r_count_25_io_out ? io_r_138_b : _GEN_10317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10319 = 9'h8b == r_count_25_io_out ? io_r_139_b : _GEN_10318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10320 = 9'h8c == r_count_25_io_out ? io_r_140_b : _GEN_10319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10321 = 9'h8d == r_count_25_io_out ? io_r_141_b : _GEN_10320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10322 = 9'h8e == r_count_25_io_out ? io_r_142_b : _GEN_10321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10323 = 9'h8f == r_count_25_io_out ? io_r_143_b : _GEN_10322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10324 = 9'h90 == r_count_25_io_out ? io_r_144_b : _GEN_10323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10325 = 9'h91 == r_count_25_io_out ? io_r_145_b : _GEN_10324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10326 = 9'h92 == r_count_25_io_out ? io_r_146_b : _GEN_10325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10327 = 9'h93 == r_count_25_io_out ? io_r_147_b : _GEN_10326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10328 = 9'h94 == r_count_25_io_out ? io_r_148_b : _GEN_10327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10329 = 9'h95 == r_count_25_io_out ? io_r_149_b : _GEN_10328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10330 = 9'h96 == r_count_25_io_out ? io_r_150_b : _GEN_10329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10331 = 9'h97 == r_count_25_io_out ? io_r_151_b : _GEN_10330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10332 = 9'h98 == r_count_25_io_out ? io_r_152_b : _GEN_10331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10333 = 9'h99 == r_count_25_io_out ? io_r_153_b : _GEN_10332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10334 = 9'h9a == r_count_25_io_out ? io_r_154_b : _GEN_10333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10335 = 9'h9b == r_count_25_io_out ? io_r_155_b : _GEN_10334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10336 = 9'h9c == r_count_25_io_out ? io_r_156_b : _GEN_10335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10337 = 9'h9d == r_count_25_io_out ? io_r_157_b : _GEN_10336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10338 = 9'h9e == r_count_25_io_out ? io_r_158_b : _GEN_10337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10339 = 9'h9f == r_count_25_io_out ? io_r_159_b : _GEN_10338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10340 = 9'ha0 == r_count_25_io_out ? io_r_160_b : _GEN_10339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10341 = 9'ha1 == r_count_25_io_out ? io_r_161_b : _GEN_10340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10342 = 9'ha2 == r_count_25_io_out ? io_r_162_b : _GEN_10341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10343 = 9'ha3 == r_count_25_io_out ? io_r_163_b : _GEN_10342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10344 = 9'ha4 == r_count_25_io_out ? io_r_164_b : _GEN_10343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10345 = 9'ha5 == r_count_25_io_out ? io_r_165_b : _GEN_10344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10346 = 9'ha6 == r_count_25_io_out ? io_r_166_b : _GEN_10345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10347 = 9'ha7 == r_count_25_io_out ? io_r_167_b : _GEN_10346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10348 = 9'ha8 == r_count_25_io_out ? io_r_168_b : _GEN_10347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10349 = 9'ha9 == r_count_25_io_out ? io_r_169_b : _GEN_10348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10350 = 9'haa == r_count_25_io_out ? io_r_170_b : _GEN_10349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10351 = 9'hab == r_count_25_io_out ? io_r_171_b : _GEN_10350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10352 = 9'hac == r_count_25_io_out ? io_r_172_b : _GEN_10351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10353 = 9'had == r_count_25_io_out ? io_r_173_b : _GEN_10352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10354 = 9'hae == r_count_25_io_out ? io_r_174_b : _GEN_10353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10355 = 9'haf == r_count_25_io_out ? io_r_175_b : _GEN_10354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10356 = 9'hb0 == r_count_25_io_out ? io_r_176_b : _GEN_10355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10357 = 9'hb1 == r_count_25_io_out ? io_r_177_b : _GEN_10356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10358 = 9'hb2 == r_count_25_io_out ? io_r_178_b : _GEN_10357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10359 = 9'hb3 == r_count_25_io_out ? io_r_179_b : _GEN_10358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10360 = 9'hb4 == r_count_25_io_out ? io_r_180_b : _GEN_10359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10361 = 9'hb5 == r_count_25_io_out ? io_r_181_b : _GEN_10360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10362 = 9'hb6 == r_count_25_io_out ? io_r_182_b : _GEN_10361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10363 = 9'hb7 == r_count_25_io_out ? io_r_183_b : _GEN_10362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10364 = 9'hb8 == r_count_25_io_out ? io_r_184_b : _GEN_10363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10365 = 9'hb9 == r_count_25_io_out ? io_r_185_b : _GEN_10364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10366 = 9'hba == r_count_25_io_out ? io_r_186_b : _GEN_10365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10367 = 9'hbb == r_count_25_io_out ? io_r_187_b : _GEN_10366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10368 = 9'hbc == r_count_25_io_out ? io_r_188_b : _GEN_10367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10369 = 9'hbd == r_count_25_io_out ? io_r_189_b : _GEN_10368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10370 = 9'hbe == r_count_25_io_out ? io_r_190_b : _GEN_10369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10371 = 9'hbf == r_count_25_io_out ? io_r_191_b : _GEN_10370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10372 = 9'hc0 == r_count_25_io_out ? io_r_192_b : _GEN_10371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10373 = 9'hc1 == r_count_25_io_out ? io_r_193_b : _GEN_10372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10374 = 9'hc2 == r_count_25_io_out ? io_r_194_b : _GEN_10373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10375 = 9'hc3 == r_count_25_io_out ? io_r_195_b : _GEN_10374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10376 = 9'hc4 == r_count_25_io_out ? io_r_196_b : _GEN_10375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10377 = 9'hc5 == r_count_25_io_out ? io_r_197_b : _GEN_10376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10378 = 9'hc6 == r_count_25_io_out ? io_r_198_b : _GEN_10377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10379 = 9'hc7 == r_count_25_io_out ? io_r_199_b : _GEN_10378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10380 = 9'hc8 == r_count_25_io_out ? io_r_200_b : _GEN_10379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10381 = 9'hc9 == r_count_25_io_out ? io_r_201_b : _GEN_10380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10382 = 9'hca == r_count_25_io_out ? io_r_202_b : _GEN_10381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10383 = 9'hcb == r_count_25_io_out ? io_r_203_b : _GEN_10382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10384 = 9'hcc == r_count_25_io_out ? io_r_204_b : _GEN_10383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10385 = 9'hcd == r_count_25_io_out ? io_r_205_b : _GEN_10384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10386 = 9'hce == r_count_25_io_out ? io_r_206_b : _GEN_10385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10387 = 9'hcf == r_count_25_io_out ? io_r_207_b : _GEN_10386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10388 = 9'hd0 == r_count_25_io_out ? io_r_208_b : _GEN_10387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10389 = 9'hd1 == r_count_25_io_out ? io_r_209_b : _GEN_10388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10390 = 9'hd2 == r_count_25_io_out ? io_r_210_b : _GEN_10389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10391 = 9'hd3 == r_count_25_io_out ? io_r_211_b : _GEN_10390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10392 = 9'hd4 == r_count_25_io_out ? io_r_212_b : _GEN_10391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10393 = 9'hd5 == r_count_25_io_out ? io_r_213_b : _GEN_10392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10394 = 9'hd6 == r_count_25_io_out ? io_r_214_b : _GEN_10393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10395 = 9'hd7 == r_count_25_io_out ? io_r_215_b : _GEN_10394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10396 = 9'hd8 == r_count_25_io_out ? io_r_216_b : _GEN_10395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10397 = 9'hd9 == r_count_25_io_out ? io_r_217_b : _GEN_10396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10398 = 9'hda == r_count_25_io_out ? io_r_218_b : _GEN_10397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10399 = 9'hdb == r_count_25_io_out ? io_r_219_b : _GEN_10398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10400 = 9'hdc == r_count_25_io_out ? io_r_220_b : _GEN_10399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10401 = 9'hdd == r_count_25_io_out ? io_r_221_b : _GEN_10400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10402 = 9'hde == r_count_25_io_out ? io_r_222_b : _GEN_10401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10403 = 9'hdf == r_count_25_io_out ? io_r_223_b : _GEN_10402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10404 = 9'he0 == r_count_25_io_out ? io_r_224_b : _GEN_10403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10405 = 9'he1 == r_count_25_io_out ? io_r_225_b : _GEN_10404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10406 = 9'he2 == r_count_25_io_out ? io_r_226_b : _GEN_10405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10407 = 9'he3 == r_count_25_io_out ? io_r_227_b : _GEN_10406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10408 = 9'he4 == r_count_25_io_out ? io_r_228_b : _GEN_10407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10409 = 9'he5 == r_count_25_io_out ? io_r_229_b : _GEN_10408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10410 = 9'he6 == r_count_25_io_out ? io_r_230_b : _GEN_10409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10411 = 9'he7 == r_count_25_io_out ? io_r_231_b : _GEN_10410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10412 = 9'he8 == r_count_25_io_out ? io_r_232_b : _GEN_10411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10413 = 9'he9 == r_count_25_io_out ? io_r_233_b : _GEN_10412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10414 = 9'hea == r_count_25_io_out ? io_r_234_b : _GEN_10413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10415 = 9'heb == r_count_25_io_out ? io_r_235_b : _GEN_10414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10416 = 9'hec == r_count_25_io_out ? io_r_236_b : _GEN_10415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10417 = 9'hed == r_count_25_io_out ? io_r_237_b : _GEN_10416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10418 = 9'hee == r_count_25_io_out ? io_r_238_b : _GEN_10417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10419 = 9'hef == r_count_25_io_out ? io_r_239_b : _GEN_10418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10420 = 9'hf0 == r_count_25_io_out ? io_r_240_b : _GEN_10419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10421 = 9'hf1 == r_count_25_io_out ? io_r_241_b : _GEN_10420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10422 = 9'hf2 == r_count_25_io_out ? io_r_242_b : _GEN_10421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10423 = 9'hf3 == r_count_25_io_out ? io_r_243_b : _GEN_10422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10424 = 9'hf4 == r_count_25_io_out ? io_r_244_b : _GEN_10423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10425 = 9'hf5 == r_count_25_io_out ? io_r_245_b : _GEN_10424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10426 = 9'hf6 == r_count_25_io_out ? io_r_246_b : _GEN_10425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10427 = 9'hf7 == r_count_25_io_out ? io_r_247_b : _GEN_10426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10428 = 9'hf8 == r_count_25_io_out ? io_r_248_b : _GEN_10427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10429 = 9'hf9 == r_count_25_io_out ? io_r_249_b : _GEN_10428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10430 = 9'hfa == r_count_25_io_out ? io_r_250_b : _GEN_10429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10431 = 9'hfb == r_count_25_io_out ? io_r_251_b : _GEN_10430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10432 = 9'hfc == r_count_25_io_out ? io_r_252_b : _GEN_10431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10433 = 9'hfd == r_count_25_io_out ? io_r_253_b : _GEN_10432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10434 = 9'hfe == r_count_25_io_out ? io_r_254_b : _GEN_10433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10435 = 9'hff == r_count_25_io_out ? io_r_255_b : _GEN_10434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10436 = 9'h100 == r_count_25_io_out ? io_r_256_b : _GEN_10435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10437 = 9'h101 == r_count_25_io_out ? io_r_257_b : _GEN_10436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10438 = 9'h102 == r_count_25_io_out ? io_r_258_b : _GEN_10437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10439 = 9'h103 == r_count_25_io_out ? io_r_259_b : _GEN_10438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10440 = 9'h104 == r_count_25_io_out ? io_r_260_b : _GEN_10439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10441 = 9'h105 == r_count_25_io_out ? io_r_261_b : _GEN_10440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10442 = 9'h106 == r_count_25_io_out ? io_r_262_b : _GEN_10441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10443 = 9'h107 == r_count_25_io_out ? io_r_263_b : _GEN_10442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10444 = 9'h108 == r_count_25_io_out ? io_r_264_b : _GEN_10443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10445 = 9'h109 == r_count_25_io_out ? io_r_265_b : _GEN_10444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10446 = 9'h10a == r_count_25_io_out ? io_r_266_b : _GEN_10445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10447 = 9'h10b == r_count_25_io_out ? io_r_267_b : _GEN_10446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10448 = 9'h10c == r_count_25_io_out ? io_r_268_b : _GEN_10447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10449 = 9'h10d == r_count_25_io_out ? io_r_269_b : _GEN_10448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10450 = 9'h10e == r_count_25_io_out ? io_r_270_b : _GEN_10449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10451 = 9'h10f == r_count_25_io_out ? io_r_271_b : _GEN_10450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10452 = 9'h110 == r_count_25_io_out ? io_r_272_b : _GEN_10451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10453 = 9'h111 == r_count_25_io_out ? io_r_273_b : _GEN_10452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10454 = 9'h112 == r_count_25_io_out ? io_r_274_b : _GEN_10453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10455 = 9'h113 == r_count_25_io_out ? io_r_275_b : _GEN_10454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10456 = 9'h114 == r_count_25_io_out ? io_r_276_b : _GEN_10455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10457 = 9'h115 == r_count_25_io_out ? io_r_277_b : _GEN_10456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10458 = 9'h116 == r_count_25_io_out ? io_r_278_b : _GEN_10457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10459 = 9'h117 == r_count_25_io_out ? io_r_279_b : _GEN_10458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10460 = 9'h118 == r_count_25_io_out ? io_r_280_b : _GEN_10459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10461 = 9'h119 == r_count_25_io_out ? io_r_281_b : _GEN_10460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10462 = 9'h11a == r_count_25_io_out ? io_r_282_b : _GEN_10461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10463 = 9'h11b == r_count_25_io_out ? io_r_283_b : _GEN_10462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10464 = 9'h11c == r_count_25_io_out ? io_r_284_b : _GEN_10463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10465 = 9'h11d == r_count_25_io_out ? io_r_285_b : _GEN_10464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10466 = 9'h11e == r_count_25_io_out ? io_r_286_b : _GEN_10465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10467 = 9'h11f == r_count_25_io_out ? io_r_287_b : _GEN_10466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10468 = 9'h120 == r_count_25_io_out ? io_r_288_b : _GEN_10467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10469 = 9'h121 == r_count_25_io_out ? io_r_289_b : _GEN_10468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10470 = 9'h122 == r_count_25_io_out ? io_r_290_b : _GEN_10469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10471 = 9'h123 == r_count_25_io_out ? io_r_291_b : _GEN_10470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10472 = 9'h124 == r_count_25_io_out ? io_r_292_b : _GEN_10471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10473 = 9'h125 == r_count_25_io_out ? io_r_293_b : _GEN_10472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10474 = 9'h126 == r_count_25_io_out ? io_r_294_b : _GEN_10473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10475 = 9'h127 == r_count_25_io_out ? io_r_295_b : _GEN_10474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10476 = 9'h128 == r_count_25_io_out ? io_r_296_b : _GEN_10475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10477 = 9'h129 == r_count_25_io_out ? io_r_297_b : _GEN_10476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10478 = 9'h12a == r_count_25_io_out ? io_r_298_b : _GEN_10477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10479 = 9'h12b == r_count_25_io_out ? io_r_299_b : _GEN_10478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10480 = 9'h12c == r_count_25_io_out ? io_r_300_b : _GEN_10479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10481 = 9'h12d == r_count_25_io_out ? io_r_301_b : _GEN_10480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10482 = 9'h12e == r_count_25_io_out ? io_r_302_b : _GEN_10481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10483 = 9'h12f == r_count_25_io_out ? io_r_303_b : _GEN_10482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10484 = 9'h130 == r_count_25_io_out ? io_r_304_b : _GEN_10483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10485 = 9'h131 == r_count_25_io_out ? io_r_305_b : _GEN_10484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10486 = 9'h132 == r_count_25_io_out ? io_r_306_b : _GEN_10485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10487 = 9'h133 == r_count_25_io_out ? io_r_307_b : _GEN_10486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10488 = 9'h134 == r_count_25_io_out ? io_r_308_b : _GEN_10487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10489 = 9'h135 == r_count_25_io_out ? io_r_309_b : _GEN_10488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10490 = 9'h136 == r_count_25_io_out ? io_r_310_b : _GEN_10489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10491 = 9'h137 == r_count_25_io_out ? io_r_311_b : _GEN_10490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10492 = 9'h138 == r_count_25_io_out ? io_r_312_b : _GEN_10491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10493 = 9'h139 == r_count_25_io_out ? io_r_313_b : _GEN_10492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10494 = 9'h13a == r_count_25_io_out ? io_r_314_b : _GEN_10493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10495 = 9'h13b == r_count_25_io_out ? io_r_315_b : _GEN_10494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10496 = 9'h13c == r_count_25_io_out ? io_r_316_b : _GEN_10495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10497 = 9'h13d == r_count_25_io_out ? io_r_317_b : _GEN_10496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10498 = 9'h13e == r_count_25_io_out ? io_r_318_b : _GEN_10497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10499 = 9'h13f == r_count_25_io_out ? io_r_319_b : _GEN_10498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10500 = 9'h140 == r_count_25_io_out ? io_r_320_b : _GEN_10499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10501 = 9'h141 == r_count_25_io_out ? io_r_321_b : _GEN_10500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10502 = 9'h142 == r_count_25_io_out ? io_r_322_b : _GEN_10501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10503 = 9'h143 == r_count_25_io_out ? io_r_323_b : _GEN_10502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10504 = 9'h144 == r_count_25_io_out ? io_r_324_b : _GEN_10503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10505 = 9'h145 == r_count_25_io_out ? io_r_325_b : _GEN_10504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10506 = 9'h146 == r_count_25_io_out ? io_r_326_b : _GEN_10505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10507 = 9'h147 == r_count_25_io_out ? io_r_327_b : _GEN_10506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10508 = 9'h148 == r_count_25_io_out ? io_r_328_b : _GEN_10507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10509 = 9'h149 == r_count_25_io_out ? io_r_329_b : _GEN_10508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10510 = 9'h14a == r_count_25_io_out ? io_r_330_b : _GEN_10509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10511 = 9'h14b == r_count_25_io_out ? io_r_331_b : _GEN_10510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10512 = 9'h14c == r_count_25_io_out ? io_r_332_b : _GEN_10511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10513 = 9'h14d == r_count_25_io_out ? io_r_333_b : _GEN_10512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10514 = 9'h14e == r_count_25_io_out ? io_r_334_b : _GEN_10513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10515 = 9'h14f == r_count_25_io_out ? io_r_335_b : _GEN_10514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10516 = 9'h150 == r_count_25_io_out ? io_r_336_b : _GEN_10515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10517 = 9'h151 == r_count_25_io_out ? io_r_337_b : _GEN_10516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10518 = 9'h152 == r_count_25_io_out ? io_r_338_b : _GEN_10517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10519 = 9'h153 == r_count_25_io_out ? io_r_339_b : _GEN_10518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10520 = 9'h154 == r_count_25_io_out ? io_r_340_b : _GEN_10519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10521 = 9'h155 == r_count_25_io_out ? io_r_341_b : _GEN_10520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10522 = 9'h156 == r_count_25_io_out ? io_r_342_b : _GEN_10521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10523 = 9'h157 == r_count_25_io_out ? io_r_343_b : _GEN_10522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10524 = 9'h158 == r_count_25_io_out ? io_r_344_b : _GEN_10523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10525 = 9'h159 == r_count_25_io_out ? io_r_345_b : _GEN_10524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10526 = 9'h15a == r_count_25_io_out ? io_r_346_b : _GEN_10525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10527 = 9'h15b == r_count_25_io_out ? io_r_347_b : _GEN_10526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10528 = 9'h15c == r_count_25_io_out ? io_r_348_b : _GEN_10527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10529 = 9'h15d == r_count_25_io_out ? io_r_349_b : _GEN_10528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10530 = 9'h15e == r_count_25_io_out ? io_r_350_b : _GEN_10529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10531 = 9'h15f == r_count_25_io_out ? io_r_351_b : _GEN_10530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10532 = 9'h160 == r_count_25_io_out ? io_r_352_b : _GEN_10531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10533 = 9'h161 == r_count_25_io_out ? io_r_353_b : _GEN_10532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10534 = 9'h162 == r_count_25_io_out ? io_r_354_b : _GEN_10533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10535 = 9'h163 == r_count_25_io_out ? io_r_355_b : _GEN_10534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10536 = 9'h164 == r_count_25_io_out ? io_r_356_b : _GEN_10535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10537 = 9'h165 == r_count_25_io_out ? io_r_357_b : _GEN_10536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10538 = 9'h166 == r_count_25_io_out ? io_r_358_b : _GEN_10537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10539 = 9'h167 == r_count_25_io_out ? io_r_359_b : _GEN_10538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10540 = 9'h168 == r_count_25_io_out ? io_r_360_b : _GEN_10539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10541 = 9'h169 == r_count_25_io_out ? io_r_361_b : _GEN_10540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10542 = 9'h16a == r_count_25_io_out ? io_r_362_b : _GEN_10541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10543 = 9'h16b == r_count_25_io_out ? io_r_363_b : _GEN_10542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10544 = 9'h16c == r_count_25_io_out ? io_r_364_b : _GEN_10543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10545 = 9'h16d == r_count_25_io_out ? io_r_365_b : _GEN_10544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10546 = 9'h16e == r_count_25_io_out ? io_r_366_b : _GEN_10545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10547 = 9'h16f == r_count_25_io_out ? io_r_367_b : _GEN_10546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10548 = 9'h170 == r_count_25_io_out ? io_r_368_b : _GEN_10547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10549 = 9'h171 == r_count_25_io_out ? io_r_369_b : _GEN_10548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10550 = 9'h172 == r_count_25_io_out ? io_r_370_b : _GEN_10549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10551 = 9'h173 == r_count_25_io_out ? io_r_371_b : _GEN_10550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10552 = 9'h174 == r_count_25_io_out ? io_r_372_b : _GEN_10551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10553 = 9'h175 == r_count_25_io_out ? io_r_373_b : _GEN_10552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10554 = 9'h176 == r_count_25_io_out ? io_r_374_b : _GEN_10553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10555 = 9'h177 == r_count_25_io_out ? io_r_375_b : _GEN_10554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10556 = 9'h178 == r_count_25_io_out ? io_r_376_b : _GEN_10555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10557 = 9'h179 == r_count_25_io_out ? io_r_377_b : _GEN_10556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10558 = 9'h17a == r_count_25_io_out ? io_r_378_b : _GEN_10557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10559 = 9'h17b == r_count_25_io_out ? io_r_379_b : _GEN_10558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10560 = 9'h17c == r_count_25_io_out ? io_r_380_b : _GEN_10559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10561 = 9'h17d == r_count_25_io_out ? io_r_381_b : _GEN_10560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10562 = 9'h17e == r_count_25_io_out ? io_r_382_b : _GEN_10561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10563 = 9'h17f == r_count_25_io_out ? io_r_383_b : _GEN_10562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10564 = 9'h180 == r_count_25_io_out ? io_r_384_b : _GEN_10563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10565 = 9'h181 == r_count_25_io_out ? io_r_385_b : _GEN_10564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10566 = 9'h182 == r_count_25_io_out ? io_r_386_b : _GEN_10565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10567 = 9'h183 == r_count_25_io_out ? io_r_387_b : _GEN_10566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10568 = 9'h184 == r_count_25_io_out ? io_r_388_b : _GEN_10567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10569 = 9'h185 == r_count_25_io_out ? io_r_389_b : _GEN_10568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10570 = 9'h186 == r_count_25_io_out ? io_r_390_b : _GEN_10569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10571 = 9'h187 == r_count_25_io_out ? io_r_391_b : _GEN_10570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10572 = 9'h188 == r_count_25_io_out ? io_r_392_b : _GEN_10571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10573 = 9'h189 == r_count_25_io_out ? io_r_393_b : _GEN_10572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10574 = 9'h18a == r_count_25_io_out ? io_r_394_b : _GEN_10573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10575 = 9'h18b == r_count_25_io_out ? io_r_395_b : _GEN_10574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10576 = 9'h18c == r_count_25_io_out ? io_r_396_b : _GEN_10575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10577 = 9'h18d == r_count_25_io_out ? io_r_397_b : _GEN_10576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10578 = 9'h18e == r_count_25_io_out ? io_r_398_b : _GEN_10577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10581 = 9'h1 == r_count_26_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10582 = 9'h2 == r_count_26_io_out ? io_r_2_b : _GEN_10581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10583 = 9'h3 == r_count_26_io_out ? io_r_3_b : _GEN_10582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10584 = 9'h4 == r_count_26_io_out ? io_r_4_b : _GEN_10583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10585 = 9'h5 == r_count_26_io_out ? io_r_5_b : _GEN_10584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10586 = 9'h6 == r_count_26_io_out ? io_r_6_b : _GEN_10585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10587 = 9'h7 == r_count_26_io_out ? io_r_7_b : _GEN_10586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10588 = 9'h8 == r_count_26_io_out ? io_r_8_b : _GEN_10587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10589 = 9'h9 == r_count_26_io_out ? io_r_9_b : _GEN_10588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10590 = 9'ha == r_count_26_io_out ? io_r_10_b : _GEN_10589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10591 = 9'hb == r_count_26_io_out ? io_r_11_b : _GEN_10590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10592 = 9'hc == r_count_26_io_out ? io_r_12_b : _GEN_10591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10593 = 9'hd == r_count_26_io_out ? io_r_13_b : _GEN_10592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10594 = 9'he == r_count_26_io_out ? io_r_14_b : _GEN_10593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10595 = 9'hf == r_count_26_io_out ? io_r_15_b : _GEN_10594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10596 = 9'h10 == r_count_26_io_out ? io_r_16_b : _GEN_10595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10597 = 9'h11 == r_count_26_io_out ? io_r_17_b : _GEN_10596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10598 = 9'h12 == r_count_26_io_out ? io_r_18_b : _GEN_10597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10599 = 9'h13 == r_count_26_io_out ? io_r_19_b : _GEN_10598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10600 = 9'h14 == r_count_26_io_out ? io_r_20_b : _GEN_10599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10601 = 9'h15 == r_count_26_io_out ? io_r_21_b : _GEN_10600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10602 = 9'h16 == r_count_26_io_out ? io_r_22_b : _GEN_10601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10603 = 9'h17 == r_count_26_io_out ? io_r_23_b : _GEN_10602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10604 = 9'h18 == r_count_26_io_out ? io_r_24_b : _GEN_10603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10605 = 9'h19 == r_count_26_io_out ? io_r_25_b : _GEN_10604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10606 = 9'h1a == r_count_26_io_out ? io_r_26_b : _GEN_10605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10607 = 9'h1b == r_count_26_io_out ? io_r_27_b : _GEN_10606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10608 = 9'h1c == r_count_26_io_out ? io_r_28_b : _GEN_10607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10609 = 9'h1d == r_count_26_io_out ? io_r_29_b : _GEN_10608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10610 = 9'h1e == r_count_26_io_out ? io_r_30_b : _GEN_10609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10611 = 9'h1f == r_count_26_io_out ? io_r_31_b : _GEN_10610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10612 = 9'h20 == r_count_26_io_out ? io_r_32_b : _GEN_10611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10613 = 9'h21 == r_count_26_io_out ? io_r_33_b : _GEN_10612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10614 = 9'h22 == r_count_26_io_out ? io_r_34_b : _GEN_10613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10615 = 9'h23 == r_count_26_io_out ? io_r_35_b : _GEN_10614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10616 = 9'h24 == r_count_26_io_out ? io_r_36_b : _GEN_10615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10617 = 9'h25 == r_count_26_io_out ? io_r_37_b : _GEN_10616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10618 = 9'h26 == r_count_26_io_out ? io_r_38_b : _GEN_10617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10619 = 9'h27 == r_count_26_io_out ? io_r_39_b : _GEN_10618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10620 = 9'h28 == r_count_26_io_out ? io_r_40_b : _GEN_10619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10621 = 9'h29 == r_count_26_io_out ? io_r_41_b : _GEN_10620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10622 = 9'h2a == r_count_26_io_out ? io_r_42_b : _GEN_10621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10623 = 9'h2b == r_count_26_io_out ? io_r_43_b : _GEN_10622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10624 = 9'h2c == r_count_26_io_out ? io_r_44_b : _GEN_10623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10625 = 9'h2d == r_count_26_io_out ? io_r_45_b : _GEN_10624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10626 = 9'h2e == r_count_26_io_out ? io_r_46_b : _GEN_10625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10627 = 9'h2f == r_count_26_io_out ? io_r_47_b : _GEN_10626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10628 = 9'h30 == r_count_26_io_out ? io_r_48_b : _GEN_10627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10629 = 9'h31 == r_count_26_io_out ? io_r_49_b : _GEN_10628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10630 = 9'h32 == r_count_26_io_out ? io_r_50_b : _GEN_10629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10631 = 9'h33 == r_count_26_io_out ? io_r_51_b : _GEN_10630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10632 = 9'h34 == r_count_26_io_out ? io_r_52_b : _GEN_10631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10633 = 9'h35 == r_count_26_io_out ? io_r_53_b : _GEN_10632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10634 = 9'h36 == r_count_26_io_out ? io_r_54_b : _GEN_10633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10635 = 9'h37 == r_count_26_io_out ? io_r_55_b : _GEN_10634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10636 = 9'h38 == r_count_26_io_out ? io_r_56_b : _GEN_10635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10637 = 9'h39 == r_count_26_io_out ? io_r_57_b : _GEN_10636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10638 = 9'h3a == r_count_26_io_out ? io_r_58_b : _GEN_10637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10639 = 9'h3b == r_count_26_io_out ? io_r_59_b : _GEN_10638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10640 = 9'h3c == r_count_26_io_out ? io_r_60_b : _GEN_10639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10641 = 9'h3d == r_count_26_io_out ? io_r_61_b : _GEN_10640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10642 = 9'h3e == r_count_26_io_out ? io_r_62_b : _GEN_10641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10643 = 9'h3f == r_count_26_io_out ? io_r_63_b : _GEN_10642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10644 = 9'h40 == r_count_26_io_out ? io_r_64_b : _GEN_10643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10645 = 9'h41 == r_count_26_io_out ? io_r_65_b : _GEN_10644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10646 = 9'h42 == r_count_26_io_out ? io_r_66_b : _GEN_10645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10647 = 9'h43 == r_count_26_io_out ? io_r_67_b : _GEN_10646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10648 = 9'h44 == r_count_26_io_out ? io_r_68_b : _GEN_10647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10649 = 9'h45 == r_count_26_io_out ? io_r_69_b : _GEN_10648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10650 = 9'h46 == r_count_26_io_out ? io_r_70_b : _GEN_10649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10651 = 9'h47 == r_count_26_io_out ? io_r_71_b : _GEN_10650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10652 = 9'h48 == r_count_26_io_out ? io_r_72_b : _GEN_10651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10653 = 9'h49 == r_count_26_io_out ? io_r_73_b : _GEN_10652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10654 = 9'h4a == r_count_26_io_out ? io_r_74_b : _GEN_10653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10655 = 9'h4b == r_count_26_io_out ? io_r_75_b : _GEN_10654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10656 = 9'h4c == r_count_26_io_out ? io_r_76_b : _GEN_10655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10657 = 9'h4d == r_count_26_io_out ? io_r_77_b : _GEN_10656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10658 = 9'h4e == r_count_26_io_out ? io_r_78_b : _GEN_10657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10659 = 9'h4f == r_count_26_io_out ? io_r_79_b : _GEN_10658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10660 = 9'h50 == r_count_26_io_out ? io_r_80_b : _GEN_10659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10661 = 9'h51 == r_count_26_io_out ? io_r_81_b : _GEN_10660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10662 = 9'h52 == r_count_26_io_out ? io_r_82_b : _GEN_10661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10663 = 9'h53 == r_count_26_io_out ? io_r_83_b : _GEN_10662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10664 = 9'h54 == r_count_26_io_out ? io_r_84_b : _GEN_10663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10665 = 9'h55 == r_count_26_io_out ? io_r_85_b : _GEN_10664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10666 = 9'h56 == r_count_26_io_out ? io_r_86_b : _GEN_10665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10667 = 9'h57 == r_count_26_io_out ? io_r_87_b : _GEN_10666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10668 = 9'h58 == r_count_26_io_out ? io_r_88_b : _GEN_10667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10669 = 9'h59 == r_count_26_io_out ? io_r_89_b : _GEN_10668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10670 = 9'h5a == r_count_26_io_out ? io_r_90_b : _GEN_10669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10671 = 9'h5b == r_count_26_io_out ? io_r_91_b : _GEN_10670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10672 = 9'h5c == r_count_26_io_out ? io_r_92_b : _GEN_10671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10673 = 9'h5d == r_count_26_io_out ? io_r_93_b : _GEN_10672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10674 = 9'h5e == r_count_26_io_out ? io_r_94_b : _GEN_10673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10675 = 9'h5f == r_count_26_io_out ? io_r_95_b : _GEN_10674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10676 = 9'h60 == r_count_26_io_out ? io_r_96_b : _GEN_10675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10677 = 9'h61 == r_count_26_io_out ? io_r_97_b : _GEN_10676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10678 = 9'h62 == r_count_26_io_out ? io_r_98_b : _GEN_10677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10679 = 9'h63 == r_count_26_io_out ? io_r_99_b : _GEN_10678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10680 = 9'h64 == r_count_26_io_out ? io_r_100_b : _GEN_10679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10681 = 9'h65 == r_count_26_io_out ? io_r_101_b : _GEN_10680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10682 = 9'h66 == r_count_26_io_out ? io_r_102_b : _GEN_10681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10683 = 9'h67 == r_count_26_io_out ? io_r_103_b : _GEN_10682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10684 = 9'h68 == r_count_26_io_out ? io_r_104_b : _GEN_10683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10685 = 9'h69 == r_count_26_io_out ? io_r_105_b : _GEN_10684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10686 = 9'h6a == r_count_26_io_out ? io_r_106_b : _GEN_10685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10687 = 9'h6b == r_count_26_io_out ? io_r_107_b : _GEN_10686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10688 = 9'h6c == r_count_26_io_out ? io_r_108_b : _GEN_10687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10689 = 9'h6d == r_count_26_io_out ? io_r_109_b : _GEN_10688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10690 = 9'h6e == r_count_26_io_out ? io_r_110_b : _GEN_10689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10691 = 9'h6f == r_count_26_io_out ? io_r_111_b : _GEN_10690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10692 = 9'h70 == r_count_26_io_out ? io_r_112_b : _GEN_10691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10693 = 9'h71 == r_count_26_io_out ? io_r_113_b : _GEN_10692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10694 = 9'h72 == r_count_26_io_out ? io_r_114_b : _GEN_10693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10695 = 9'h73 == r_count_26_io_out ? io_r_115_b : _GEN_10694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10696 = 9'h74 == r_count_26_io_out ? io_r_116_b : _GEN_10695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10697 = 9'h75 == r_count_26_io_out ? io_r_117_b : _GEN_10696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10698 = 9'h76 == r_count_26_io_out ? io_r_118_b : _GEN_10697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10699 = 9'h77 == r_count_26_io_out ? io_r_119_b : _GEN_10698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10700 = 9'h78 == r_count_26_io_out ? io_r_120_b : _GEN_10699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10701 = 9'h79 == r_count_26_io_out ? io_r_121_b : _GEN_10700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10702 = 9'h7a == r_count_26_io_out ? io_r_122_b : _GEN_10701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10703 = 9'h7b == r_count_26_io_out ? io_r_123_b : _GEN_10702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10704 = 9'h7c == r_count_26_io_out ? io_r_124_b : _GEN_10703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10705 = 9'h7d == r_count_26_io_out ? io_r_125_b : _GEN_10704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10706 = 9'h7e == r_count_26_io_out ? io_r_126_b : _GEN_10705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10707 = 9'h7f == r_count_26_io_out ? io_r_127_b : _GEN_10706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10708 = 9'h80 == r_count_26_io_out ? io_r_128_b : _GEN_10707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10709 = 9'h81 == r_count_26_io_out ? io_r_129_b : _GEN_10708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10710 = 9'h82 == r_count_26_io_out ? io_r_130_b : _GEN_10709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10711 = 9'h83 == r_count_26_io_out ? io_r_131_b : _GEN_10710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10712 = 9'h84 == r_count_26_io_out ? io_r_132_b : _GEN_10711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10713 = 9'h85 == r_count_26_io_out ? io_r_133_b : _GEN_10712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10714 = 9'h86 == r_count_26_io_out ? io_r_134_b : _GEN_10713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10715 = 9'h87 == r_count_26_io_out ? io_r_135_b : _GEN_10714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10716 = 9'h88 == r_count_26_io_out ? io_r_136_b : _GEN_10715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10717 = 9'h89 == r_count_26_io_out ? io_r_137_b : _GEN_10716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10718 = 9'h8a == r_count_26_io_out ? io_r_138_b : _GEN_10717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10719 = 9'h8b == r_count_26_io_out ? io_r_139_b : _GEN_10718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10720 = 9'h8c == r_count_26_io_out ? io_r_140_b : _GEN_10719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10721 = 9'h8d == r_count_26_io_out ? io_r_141_b : _GEN_10720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10722 = 9'h8e == r_count_26_io_out ? io_r_142_b : _GEN_10721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10723 = 9'h8f == r_count_26_io_out ? io_r_143_b : _GEN_10722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10724 = 9'h90 == r_count_26_io_out ? io_r_144_b : _GEN_10723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10725 = 9'h91 == r_count_26_io_out ? io_r_145_b : _GEN_10724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10726 = 9'h92 == r_count_26_io_out ? io_r_146_b : _GEN_10725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10727 = 9'h93 == r_count_26_io_out ? io_r_147_b : _GEN_10726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10728 = 9'h94 == r_count_26_io_out ? io_r_148_b : _GEN_10727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10729 = 9'h95 == r_count_26_io_out ? io_r_149_b : _GEN_10728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10730 = 9'h96 == r_count_26_io_out ? io_r_150_b : _GEN_10729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10731 = 9'h97 == r_count_26_io_out ? io_r_151_b : _GEN_10730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10732 = 9'h98 == r_count_26_io_out ? io_r_152_b : _GEN_10731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10733 = 9'h99 == r_count_26_io_out ? io_r_153_b : _GEN_10732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10734 = 9'h9a == r_count_26_io_out ? io_r_154_b : _GEN_10733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10735 = 9'h9b == r_count_26_io_out ? io_r_155_b : _GEN_10734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10736 = 9'h9c == r_count_26_io_out ? io_r_156_b : _GEN_10735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10737 = 9'h9d == r_count_26_io_out ? io_r_157_b : _GEN_10736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10738 = 9'h9e == r_count_26_io_out ? io_r_158_b : _GEN_10737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10739 = 9'h9f == r_count_26_io_out ? io_r_159_b : _GEN_10738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10740 = 9'ha0 == r_count_26_io_out ? io_r_160_b : _GEN_10739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10741 = 9'ha1 == r_count_26_io_out ? io_r_161_b : _GEN_10740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10742 = 9'ha2 == r_count_26_io_out ? io_r_162_b : _GEN_10741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10743 = 9'ha3 == r_count_26_io_out ? io_r_163_b : _GEN_10742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10744 = 9'ha4 == r_count_26_io_out ? io_r_164_b : _GEN_10743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10745 = 9'ha5 == r_count_26_io_out ? io_r_165_b : _GEN_10744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10746 = 9'ha6 == r_count_26_io_out ? io_r_166_b : _GEN_10745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10747 = 9'ha7 == r_count_26_io_out ? io_r_167_b : _GEN_10746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10748 = 9'ha8 == r_count_26_io_out ? io_r_168_b : _GEN_10747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10749 = 9'ha9 == r_count_26_io_out ? io_r_169_b : _GEN_10748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10750 = 9'haa == r_count_26_io_out ? io_r_170_b : _GEN_10749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10751 = 9'hab == r_count_26_io_out ? io_r_171_b : _GEN_10750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10752 = 9'hac == r_count_26_io_out ? io_r_172_b : _GEN_10751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10753 = 9'had == r_count_26_io_out ? io_r_173_b : _GEN_10752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10754 = 9'hae == r_count_26_io_out ? io_r_174_b : _GEN_10753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10755 = 9'haf == r_count_26_io_out ? io_r_175_b : _GEN_10754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10756 = 9'hb0 == r_count_26_io_out ? io_r_176_b : _GEN_10755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10757 = 9'hb1 == r_count_26_io_out ? io_r_177_b : _GEN_10756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10758 = 9'hb2 == r_count_26_io_out ? io_r_178_b : _GEN_10757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10759 = 9'hb3 == r_count_26_io_out ? io_r_179_b : _GEN_10758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10760 = 9'hb4 == r_count_26_io_out ? io_r_180_b : _GEN_10759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10761 = 9'hb5 == r_count_26_io_out ? io_r_181_b : _GEN_10760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10762 = 9'hb6 == r_count_26_io_out ? io_r_182_b : _GEN_10761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10763 = 9'hb7 == r_count_26_io_out ? io_r_183_b : _GEN_10762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10764 = 9'hb8 == r_count_26_io_out ? io_r_184_b : _GEN_10763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10765 = 9'hb9 == r_count_26_io_out ? io_r_185_b : _GEN_10764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10766 = 9'hba == r_count_26_io_out ? io_r_186_b : _GEN_10765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10767 = 9'hbb == r_count_26_io_out ? io_r_187_b : _GEN_10766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10768 = 9'hbc == r_count_26_io_out ? io_r_188_b : _GEN_10767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10769 = 9'hbd == r_count_26_io_out ? io_r_189_b : _GEN_10768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10770 = 9'hbe == r_count_26_io_out ? io_r_190_b : _GEN_10769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10771 = 9'hbf == r_count_26_io_out ? io_r_191_b : _GEN_10770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10772 = 9'hc0 == r_count_26_io_out ? io_r_192_b : _GEN_10771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10773 = 9'hc1 == r_count_26_io_out ? io_r_193_b : _GEN_10772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10774 = 9'hc2 == r_count_26_io_out ? io_r_194_b : _GEN_10773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10775 = 9'hc3 == r_count_26_io_out ? io_r_195_b : _GEN_10774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10776 = 9'hc4 == r_count_26_io_out ? io_r_196_b : _GEN_10775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10777 = 9'hc5 == r_count_26_io_out ? io_r_197_b : _GEN_10776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10778 = 9'hc6 == r_count_26_io_out ? io_r_198_b : _GEN_10777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10779 = 9'hc7 == r_count_26_io_out ? io_r_199_b : _GEN_10778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10780 = 9'hc8 == r_count_26_io_out ? io_r_200_b : _GEN_10779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10781 = 9'hc9 == r_count_26_io_out ? io_r_201_b : _GEN_10780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10782 = 9'hca == r_count_26_io_out ? io_r_202_b : _GEN_10781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10783 = 9'hcb == r_count_26_io_out ? io_r_203_b : _GEN_10782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10784 = 9'hcc == r_count_26_io_out ? io_r_204_b : _GEN_10783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10785 = 9'hcd == r_count_26_io_out ? io_r_205_b : _GEN_10784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10786 = 9'hce == r_count_26_io_out ? io_r_206_b : _GEN_10785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10787 = 9'hcf == r_count_26_io_out ? io_r_207_b : _GEN_10786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10788 = 9'hd0 == r_count_26_io_out ? io_r_208_b : _GEN_10787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10789 = 9'hd1 == r_count_26_io_out ? io_r_209_b : _GEN_10788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10790 = 9'hd2 == r_count_26_io_out ? io_r_210_b : _GEN_10789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10791 = 9'hd3 == r_count_26_io_out ? io_r_211_b : _GEN_10790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10792 = 9'hd4 == r_count_26_io_out ? io_r_212_b : _GEN_10791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10793 = 9'hd5 == r_count_26_io_out ? io_r_213_b : _GEN_10792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10794 = 9'hd6 == r_count_26_io_out ? io_r_214_b : _GEN_10793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10795 = 9'hd7 == r_count_26_io_out ? io_r_215_b : _GEN_10794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10796 = 9'hd8 == r_count_26_io_out ? io_r_216_b : _GEN_10795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10797 = 9'hd9 == r_count_26_io_out ? io_r_217_b : _GEN_10796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10798 = 9'hda == r_count_26_io_out ? io_r_218_b : _GEN_10797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10799 = 9'hdb == r_count_26_io_out ? io_r_219_b : _GEN_10798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10800 = 9'hdc == r_count_26_io_out ? io_r_220_b : _GEN_10799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10801 = 9'hdd == r_count_26_io_out ? io_r_221_b : _GEN_10800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10802 = 9'hde == r_count_26_io_out ? io_r_222_b : _GEN_10801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10803 = 9'hdf == r_count_26_io_out ? io_r_223_b : _GEN_10802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10804 = 9'he0 == r_count_26_io_out ? io_r_224_b : _GEN_10803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10805 = 9'he1 == r_count_26_io_out ? io_r_225_b : _GEN_10804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10806 = 9'he2 == r_count_26_io_out ? io_r_226_b : _GEN_10805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10807 = 9'he3 == r_count_26_io_out ? io_r_227_b : _GEN_10806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10808 = 9'he4 == r_count_26_io_out ? io_r_228_b : _GEN_10807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10809 = 9'he5 == r_count_26_io_out ? io_r_229_b : _GEN_10808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10810 = 9'he6 == r_count_26_io_out ? io_r_230_b : _GEN_10809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10811 = 9'he7 == r_count_26_io_out ? io_r_231_b : _GEN_10810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10812 = 9'he8 == r_count_26_io_out ? io_r_232_b : _GEN_10811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10813 = 9'he9 == r_count_26_io_out ? io_r_233_b : _GEN_10812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10814 = 9'hea == r_count_26_io_out ? io_r_234_b : _GEN_10813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10815 = 9'heb == r_count_26_io_out ? io_r_235_b : _GEN_10814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10816 = 9'hec == r_count_26_io_out ? io_r_236_b : _GEN_10815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10817 = 9'hed == r_count_26_io_out ? io_r_237_b : _GEN_10816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10818 = 9'hee == r_count_26_io_out ? io_r_238_b : _GEN_10817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10819 = 9'hef == r_count_26_io_out ? io_r_239_b : _GEN_10818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10820 = 9'hf0 == r_count_26_io_out ? io_r_240_b : _GEN_10819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10821 = 9'hf1 == r_count_26_io_out ? io_r_241_b : _GEN_10820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10822 = 9'hf2 == r_count_26_io_out ? io_r_242_b : _GEN_10821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10823 = 9'hf3 == r_count_26_io_out ? io_r_243_b : _GEN_10822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10824 = 9'hf4 == r_count_26_io_out ? io_r_244_b : _GEN_10823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10825 = 9'hf5 == r_count_26_io_out ? io_r_245_b : _GEN_10824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10826 = 9'hf6 == r_count_26_io_out ? io_r_246_b : _GEN_10825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10827 = 9'hf7 == r_count_26_io_out ? io_r_247_b : _GEN_10826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10828 = 9'hf8 == r_count_26_io_out ? io_r_248_b : _GEN_10827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10829 = 9'hf9 == r_count_26_io_out ? io_r_249_b : _GEN_10828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10830 = 9'hfa == r_count_26_io_out ? io_r_250_b : _GEN_10829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10831 = 9'hfb == r_count_26_io_out ? io_r_251_b : _GEN_10830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10832 = 9'hfc == r_count_26_io_out ? io_r_252_b : _GEN_10831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10833 = 9'hfd == r_count_26_io_out ? io_r_253_b : _GEN_10832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10834 = 9'hfe == r_count_26_io_out ? io_r_254_b : _GEN_10833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10835 = 9'hff == r_count_26_io_out ? io_r_255_b : _GEN_10834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10836 = 9'h100 == r_count_26_io_out ? io_r_256_b : _GEN_10835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10837 = 9'h101 == r_count_26_io_out ? io_r_257_b : _GEN_10836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10838 = 9'h102 == r_count_26_io_out ? io_r_258_b : _GEN_10837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10839 = 9'h103 == r_count_26_io_out ? io_r_259_b : _GEN_10838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10840 = 9'h104 == r_count_26_io_out ? io_r_260_b : _GEN_10839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10841 = 9'h105 == r_count_26_io_out ? io_r_261_b : _GEN_10840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10842 = 9'h106 == r_count_26_io_out ? io_r_262_b : _GEN_10841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10843 = 9'h107 == r_count_26_io_out ? io_r_263_b : _GEN_10842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10844 = 9'h108 == r_count_26_io_out ? io_r_264_b : _GEN_10843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10845 = 9'h109 == r_count_26_io_out ? io_r_265_b : _GEN_10844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10846 = 9'h10a == r_count_26_io_out ? io_r_266_b : _GEN_10845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10847 = 9'h10b == r_count_26_io_out ? io_r_267_b : _GEN_10846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10848 = 9'h10c == r_count_26_io_out ? io_r_268_b : _GEN_10847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10849 = 9'h10d == r_count_26_io_out ? io_r_269_b : _GEN_10848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10850 = 9'h10e == r_count_26_io_out ? io_r_270_b : _GEN_10849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10851 = 9'h10f == r_count_26_io_out ? io_r_271_b : _GEN_10850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10852 = 9'h110 == r_count_26_io_out ? io_r_272_b : _GEN_10851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10853 = 9'h111 == r_count_26_io_out ? io_r_273_b : _GEN_10852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10854 = 9'h112 == r_count_26_io_out ? io_r_274_b : _GEN_10853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10855 = 9'h113 == r_count_26_io_out ? io_r_275_b : _GEN_10854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10856 = 9'h114 == r_count_26_io_out ? io_r_276_b : _GEN_10855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10857 = 9'h115 == r_count_26_io_out ? io_r_277_b : _GEN_10856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10858 = 9'h116 == r_count_26_io_out ? io_r_278_b : _GEN_10857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10859 = 9'h117 == r_count_26_io_out ? io_r_279_b : _GEN_10858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10860 = 9'h118 == r_count_26_io_out ? io_r_280_b : _GEN_10859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10861 = 9'h119 == r_count_26_io_out ? io_r_281_b : _GEN_10860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10862 = 9'h11a == r_count_26_io_out ? io_r_282_b : _GEN_10861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10863 = 9'h11b == r_count_26_io_out ? io_r_283_b : _GEN_10862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10864 = 9'h11c == r_count_26_io_out ? io_r_284_b : _GEN_10863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10865 = 9'h11d == r_count_26_io_out ? io_r_285_b : _GEN_10864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10866 = 9'h11e == r_count_26_io_out ? io_r_286_b : _GEN_10865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10867 = 9'h11f == r_count_26_io_out ? io_r_287_b : _GEN_10866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10868 = 9'h120 == r_count_26_io_out ? io_r_288_b : _GEN_10867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10869 = 9'h121 == r_count_26_io_out ? io_r_289_b : _GEN_10868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10870 = 9'h122 == r_count_26_io_out ? io_r_290_b : _GEN_10869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10871 = 9'h123 == r_count_26_io_out ? io_r_291_b : _GEN_10870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10872 = 9'h124 == r_count_26_io_out ? io_r_292_b : _GEN_10871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10873 = 9'h125 == r_count_26_io_out ? io_r_293_b : _GEN_10872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10874 = 9'h126 == r_count_26_io_out ? io_r_294_b : _GEN_10873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10875 = 9'h127 == r_count_26_io_out ? io_r_295_b : _GEN_10874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10876 = 9'h128 == r_count_26_io_out ? io_r_296_b : _GEN_10875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10877 = 9'h129 == r_count_26_io_out ? io_r_297_b : _GEN_10876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10878 = 9'h12a == r_count_26_io_out ? io_r_298_b : _GEN_10877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10879 = 9'h12b == r_count_26_io_out ? io_r_299_b : _GEN_10878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10880 = 9'h12c == r_count_26_io_out ? io_r_300_b : _GEN_10879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10881 = 9'h12d == r_count_26_io_out ? io_r_301_b : _GEN_10880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10882 = 9'h12e == r_count_26_io_out ? io_r_302_b : _GEN_10881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10883 = 9'h12f == r_count_26_io_out ? io_r_303_b : _GEN_10882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10884 = 9'h130 == r_count_26_io_out ? io_r_304_b : _GEN_10883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10885 = 9'h131 == r_count_26_io_out ? io_r_305_b : _GEN_10884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10886 = 9'h132 == r_count_26_io_out ? io_r_306_b : _GEN_10885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10887 = 9'h133 == r_count_26_io_out ? io_r_307_b : _GEN_10886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10888 = 9'h134 == r_count_26_io_out ? io_r_308_b : _GEN_10887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10889 = 9'h135 == r_count_26_io_out ? io_r_309_b : _GEN_10888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10890 = 9'h136 == r_count_26_io_out ? io_r_310_b : _GEN_10889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10891 = 9'h137 == r_count_26_io_out ? io_r_311_b : _GEN_10890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10892 = 9'h138 == r_count_26_io_out ? io_r_312_b : _GEN_10891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10893 = 9'h139 == r_count_26_io_out ? io_r_313_b : _GEN_10892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10894 = 9'h13a == r_count_26_io_out ? io_r_314_b : _GEN_10893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10895 = 9'h13b == r_count_26_io_out ? io_r_315_b : _GEN_10894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10896 = 9'h13c == r_count_26_io_out ? io_r_316_b : _GEN_10895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10897 = 9'h13d == r_count_26_io_out ? io_r_317_b : _GEN_10896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10898 = 9'h13e == r_count_26_io_out ? io_r_318_b : _GEN_10897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10899 = 9'h13f == r_count_26_io_out ? io_r_319_b : _GEN_10898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10900 = 9'h140 == r_count_26_io_out ? io_r_320_b : _GEN_10899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10901 = 9'h141 == r_count_26_io_out ? io_r_321_b : _GEN_10900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10902 = 9'h142 == r_count_26_io_out ? io_r_322_b : _GEN_10901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10903 = 9'h143 == r_count_26_io_out ? io_r_323_b : _GEN_10902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10904 = 9'h144 == r_count_26_io_out ? io_r_324_b : _GEN_10903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10905 = 9'h145 == r_count_26_io_out ? io_r_325_b : _GEN_10904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10906 = 9'h146 == r_count_26_io_out ? io_r_326_b : _GEN_10905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10907 = 9'h147 == r_count_26_io_out ? io_r_327_b : _GEN_10906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10908 = 9'h148 == r_count_26_io_out ? io_r_328_b : _GEN_10907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10909 = 9'h149 == r_count_26_io_out ? io_r_329_b : _GEN_10908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10910 = 9'h14a == r_count_26_io_out ? io_r_330_b : _GEN_10909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10911 = 9'h14b == r_count_26_io_out ? io_r_331_b : _GEN_10910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10912 = 9'h14c == r_count_26_io_out ? io_r_332_b : _GEN_10911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10913 = 9'h14d == r_count_26_io_out ? io_r_333_b : _GEN_10912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10914 = 9'h14e == r_count_26_io_out ? io_r_334_b : _GEN_10913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10915 = 9'h14f == r_count_26_io_out ? io_r_335_b : _GEN_10914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10916 = 9'h150 == r_count_26_io_out ? io_r_336_b : _GEN_10915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10917 = 9'h151 == r_count_26_io_out ? io_r_337_b : _GEN_10916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10918 = 9'h152 == r_count_26_io_out ? io_r_338_b : _GEN_10917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10919 = 9'h153 == r_count_26_io_out ? io_r_339_b : _GEN_10918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10920 = 9'h154 == r_count_26_io_out ? io_r_340_b : _GEN_10919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10921 = 9'h155 == r_count_26_io_out ? io_r_341_b : _GEN_10920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10922 = 9'h156 == r_count_26_io_out ? io_r_342_b : _GEN_10921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10923 = 9'h157 == r_count_26_io_out ? io_r_343_b : _GEN_10922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10924 = 9'h158 == r_count_26_io_out ? io_r_344_b : _GEN_10923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10925 = 9'h159 == r_count_26_io_out ? io_r_345_b : _GEN_10924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10926 = 9'h15a == r_count_26_io_out ? io_r_346_b : _GEN_10925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10927 = 9'h15b == r_count_26_io_out ? io_r_347_b : _GEN_10926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10928 = 9'h15c == r_count_26_io_out ? io_r_348_b : _GEN_10927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10929 = 9'h15d == r_count_26_io_out ? io_r_349_b : _GEN_10928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10930 = 9'h15e == r_count_26_io_out ? io_r_350_b : _GEN_10929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10931 = 9'h15f == r_count_26_io_out ? io_r_351_b : _GEN_10930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10932 = 9'h160 == r_count_26_io_out ? io_r_352_b : _GEN_10931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10933 = 9'h161 == r_count_26_io_out ? io_r_353_b : _GEN_10932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10934 = 9'h162 == r_count_26_io_out ? io_r_354_b : _GEN_10933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10935 = 9'h163 == r_count_26_io_out ? io_r_355_b : _GEN_10934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10936 = 9'h164 == r_count_26_io_out ? io_r_356_b : _GEN_10935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10937 = 9'h165 == r_count_26_io_out ? io_r_357_b : _GEN_10936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10938 = 9'h166 == r_count_26_io_out ? io_r_358_b : _GEN_10937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10939 = 9'h167 == r_count_26_io_out ? io_r_359_b : _GEN_10938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10940 = 9'h168 == r_count_26_io_out ? io_r_360_b : _GEN_10939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10941 = 9'h169 == r_count_26_io_out ? io_r_361_b : _GEN_10940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10942 = 9'h16a == r_count_26_io_out ? io_r_362_b : _GEN_10941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10943 = 9'h16b == r_count_26_io_out ? io_r_363_b : _GEN_10942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10944 = 9'h16c == r_count_26_io_out ? io_r_364_b : _GEN_10943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10945 = 9'h16d == r_count_26_io_out ? io_r_365_b : _GEN_10944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10946 = 9'h16e == r_count_26_io_out ? io_r_366_b : _GEN_10945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10947 = 9'h16f == r_count_26_io_out ? io_r_367_b : _GEN_10946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10948 = 9'h170 == r_count_26_io_out ? io_r_368_b : _GEN_10947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10949 = 9'h171 == r_count_26_io_out ? io_r_369_b : _GEN_10948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10950 = 9'h172 == r_count_26_io_out ? io_r_370_b : _GEN_10949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10951 = 9'h173 == r_count_26_io_out ? io_r_371_b : _GEN_10950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10952 = 9'h174 == r_count_26_io_out ? io_r_372_b : _GEN_10951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10953 = 9'h175 == r_count_26_io_out ? io_r_373_b : _GEN_10952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10954 = 9'h176 == r_count_26_io_out ? io_r_374_b : _GEN_10953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10955 = 9'h177 == r_count_26_io_out ? io_r_375_b : _GEN_10954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10956 = 9'h178 == r_count_26_io_out ? io_r_376_b : _GEN_10955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10957 = 9'h179 == r_count_26_io_out ? io_r_377_b : _GEN_10956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10958 = 9'h17a == r_count_26_io_out ? io_r_378_b : _GEN_10957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10959 = 9'h17b == r_count_26_io_out ? io_r_379_b : _GEN_10958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10960 = 9'h17c == r_count_26_io_out ? io_r_380_b : _GEN_10959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10961 = 9'h17d == r_count_26_io_out ? io_r_381_b : _GEN_10960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10962 = 9'h17e == r_count_26_io_out ? io_r_382_b : _GEN_10961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10963 = 9'h17f == r_count_26_io_out ? io_r_383_b : _GEN_10962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10964 = 9'h180 == r_count_26_io_out ? io_r_384_b : _GEN_10963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10965 = 9'h181 == r_count_26_io_out ? io_r_385_b : _GEN_10964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10966 = 9'h182 == r_count_26_io_out ? io_r_386_b : _GEN_10965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10967 = 9'h183 == r_count_26_io_out ? io_r_387_b : _GEN_10966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10968 = 9'h184 == r_count_26_io_out ? io_r_388_b : _GEN_10967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10969 = 9'h185 == r_count_26_io_out ? io_r_389_b : _GEN_10968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10970 = 9'h186 == r_count_26_io_out ? io_r_390_b : _GEN_10969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10971 = 9'h187 == r_count_26_io_out ? io_r_391_b : _GEN_10970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10972 = 9'h188 == r_count_26_io_out ? io_r_392_b : _GEN_10971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10973 = 9'h189 == r_count_26_io_out ? io_r_393_b : _GEN_10972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10974 = 9'h18a == r_count_26_io_out ? io_r_394_b : _GEN_10973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10975 = 9'h18b == r_count_26_io_out ? io_r_395_b : _GEN_10974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10976 = 9'h18c == r_count_26_io_out ? io_r_396_b : _GEN_10975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10977 = 9'h18d == r_count_26_io_out ? io_r_397_b : _GEN_10976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10978 = 9'h18e == r_count_26_io_out ? io_r_398_b : _GEN_10977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10981 = 9'h1 == r_count_27_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10982 = 9'h2 == r_count_27_io_out ? io_r_2_b : _GEN_10981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10983 = 9'h3 == r_count_27_io_out ? io_r_3_b : _GEN_10982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10984 = 9'h4 == r_count_27_io_out ? io_r_4_b : _GEN_10983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10985 = 9'h5 == r_count_27_io_out ? io_r_5_b : _GEN_10984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10986 = 9'h6 == r_count_27_io_out ? io_r_6_b : _GEN_10985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10987 = 9'h7 == r_count_27_io_out ? io_r_7_b : _GEN_10986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10988 = 9'h8 == r_count_27_io_out ? io_r_8_b : _GEN_10987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10989 = 9'h9 == r_count_27_io_out ? io_r_9_b : _GEN_10988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10990 = 9'ha == r_count_27_io_out ? io_r_10_b : _GEN_10989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10991 = 9'hb == r_count_27_io_out ? io_r_11_b : _GEN_10990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10992 = 9'hc == r_count_27_io_out ? io_r_12_b : _GEN_10991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10993 = 9'hd == r_count_27_io_out ? io_r_13_b : _GEN_10992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10994 = 9'he == r_count_27_io_out ? io_r_14_b : _GEN_10993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10995 = 9'hf == r_count_27_io_out ? io_r_15_b : _GEN_10994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10996 = 9'h10 == r_count_27_io_out ? io_r_16_b : _GEN_10995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10997 = 9'h11 == r_count_27_io_out ? io_r_17_b : _GEN_10996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10998 = 9'h12 == r_count_27_io_out ? io_r_18_b : _GEN_10997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10999 = 9'h13 == r_count_27_io_out ? io_r_19_b : _GEN_10998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11000 = 9'h14 == r_count_27_io_out ? io_r_20_b : _GEN_10999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11001 = 9'h15 == r_count_27_io_out ? io_r_21_b : _GEN_11000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11002 = 9'h16 == r_count_27_io_out ? io_r_22_b : _GEN_11001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11003 = 9'h17 == r_count_27_io_out ? io_r_23_b : _GEN_11002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11004 = 9'h18 == r_count_27_io_out ? io_r_24_b : _GEN_11003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11005 = 9'h19 == r_count_27_io_out ? io_r_25_b : _GEN_11004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11006 = 9'h1a == r_count_27_io_out ? io_r_26_b : _GEN_11005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11007 = 9'h1b == r_count_27_io_out ? io_r_27_b : _GEN_11006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11008 = 9'h1c == r_count_27_io_out ? io_r_28_b : _GEN_11007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11009 = 9'h1d == r_count_27_io_out ? io_r_29_b : _GEN_11008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11010 = 9'h1e == r_count_27_io_out ? io_r_30_b : _GEN_11009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11011 = 9'h1f == r_count_27_io_out ? io_r_31_b : _GEN_11010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11012 = 9'h20 == r_count_27_io_out ? io_r_32_b : _GEN_11011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11013 = 9'h21 == r_count_27_io_out ? io_r_33_b : _GEN_11012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11014 = 9'h22 == r_count_27_io_out ? io_r_34_b : _GEN_11013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11015 = 9'h23 == r_count_27_io_out ? io_r_35_b : _GEN_11014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11016 = 9'h24 == r_count_27_io_out ? io_r_36_b : _GEN_11015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11017 = 9'h25 == r_count_27_io_out ? io_r_37_b : _GEN_11016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11018 = 9'h26 == r_count_27_io_out ? io_r_38_b : _GEN_11017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11019 = 9'h27 == r_count_27_io_out ? io_r_39_b : _GEN_11018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11020 = 9'h28 == r_count_27_io_out ? io_r_40_b : _GEN_11019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11021 = 9'h29 == r_count_27_io_out ? io_r_41_b : _GEN_11020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11022 = 9'h2a == r_count_27_io_out ? io_r_42_b : _GEN_11021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11023 = 9'h2b == r_count_27_io_out ? io_r_43_b : _GEN_11022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11024 = 9'h2c == r_count_27_io_out ? io_r_44_b : _GEN_11023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11025 = 9'h2d == r_count_27_io_out ? io_r_45_b : _GEN_11024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11026 = 9'h2e == r_count_27_io_out ? io_r_46_b : _GEN_11025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11027 = 9'h2f == r_count_27_io_out ? io_r_47_b : _GEN_11026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11028 = 9'h30 == r_count_27_io_out ? io_r_48_b : _GEN_11027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11029 = 9'h31 == r_count_27_io_out ? io_r_49_b : _GEN_11028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11030 = 9'h32 == r_count_27_io_out ? io_r_50_b : _GEN_11029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11031 = 9'h33 == r_count_27_io_out ? io_r_51_b : _GEN_11030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11032 = 9'h34 == r_count_27_io_out ? io_r_52_b : _GEN_11031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11033 = 9'h35 == r_count_27_io_out ? io_r_53_b : _GEN_11032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11034 = 9'h36 == r_count_27_io_out ? io_r_54_b : _GEN_11033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11035 = 9'h37 == r_count_27_io_out ? io_r_55_b : _GEN_11034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11036 = 9'h38 == r_count_27_io_out ? io_r_56_b : _GEN_11035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11037 = 9'h39 == r_count_27_io_out ? io_r_57_b : _GEN_11036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11038 = 9'h3a == r_count_27_io_out ? io_r_58_b : _GEN_11037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11039 = 9'h3b == r_count_27_io_out ? io_r_59_b : _GEN_11038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11040 = 9'h3c == r_count_27_io_out ? io_r_60_b : _GEN_11039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11041 = 9'h3d == r_count_27_io_out ? io_r_61_b : _GEN_11040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11042 = 9'h3e == r_count_27_io_out ? io_r_62_b : _GEN_11041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11043 = 9'h3f == r_count_27_io_out ? io_r_63_b : _GEN_11042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11044 = 9'h40 == r_count_27_io_out ? io_r_64_b : _GEN_11043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11045 = 9'h41 == r_count_27_io_out ? io_r_65_b : _GEN_11044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11046 = 9'h42 == r_count_27_io_out ? io_r_66_b : _GEN_11045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11047 = 9'h43 == r_count_27_io_out ? io_r_67_b : _GEN_11046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11048 = 9'h44 == r_count_27_io_out ? io_r_68_b : _GEN_11047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11049 = 9'h45 == r_count_27_io_out ? io_r_69_b : _GEN_11048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11050 = 9'h46 == r_count_27_io_out ? io_r_70_b : _GEN_11049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11051 = 9'h47 == r_count_27_io_out ? io_r_71_b : _GEN_11050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11052 = 9'h48 == r_count_27_io_out ? io_r_72_b : _GEN_11051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11053 = 9'h49 == r_count_27_io_out ? io_r_73_b : _GEN_11052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11054 = 9'h4a == r_count_27_io_out ? io_r_74_b : _GEN_11053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11055 = 9'h4b == r_count_27_io_out ? io_r_75_b : _GEN_11054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11056 = 9'h4c == r_count_27_io_out ? io_r_76_b : _GEN_11055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11057 = 9'h4d == r_count_27_io_out ? io_r_77_b : _GEN_11056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11058 = 9'h4e == r_count_27_io_out ? io_r_78_b : _GEN_11057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11059 = 9'h4f == r_count_27_io_out ? io_r_79_b : _GEN_11058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11060 = 9'h50 == r_count_27_io_out ? io_r_80_b : _GEN_11059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11061 = 9'h51 == r_count_27_io_out ? io_r_81_b : _GEN_11060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11062 = 9'h52 == r_count_27_io_out ? io_r_82_b : _GEN_11061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11063 = 9'h53 == r_count_27_io_out ? io_r_83_b : _GEN_11062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11064 = 9'h54 == r_count_27_io_out ? io_r_84_b : _GEN_11063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11065 = 9'h55 == r_count_27_io_out ? io_r_85_b : _GEN_11064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11066 = 9'h56 == r_count_27_io_out ? io_r_86_b : _GEN_11065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11067 = 9'h57 == r_count_27_io_out ? io_r_87_b : _GEN_11066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11068 = 9'h58 == r_count_27_io_out ? io_r_88_b : _GEN_11067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11069 = 9'h59 == r_count_27_io_out ? io_r_89_b : _GEN_11068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11070 = 9'h5a == r_count_27_io_out ? io_r_90_b : _GEN_11069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11071 = 9'h5b == r_count_27_io_out ? io_r_91_b : _GEN_11070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11072 = 9'h5c == r_count_27_io_out ? io_r_92_b : _GEN_11071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11073 = 9'h5d == r_count_27_io_out ? io_r_93_b : _GEN_11072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11074 = 9'h5e == r_count_27_io_out ? io_r_94_b : _GEN_11073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11075 = 9'h5f == r_count_27_io_out ? io_r_95_b : _GEN_11074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11076 = 9'h60 == r_count_27_io_out ? io_r_96_b : _GEN_11075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11077 = 9'h61 == r_count_27_io_out ? io_r_97_b : _GEN_11076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11078 = 9'h62 == r_count_27_io_out ? io_r_98_b : _GEN_11077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11079 = 9'h63 == r_count_27_io_out ? io_r_99_b : _GEN_11078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11080 = 9'h64 == r_count_27_io_out ? io_r_100_b : _GEN_11079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11081 = 9'h65 == r_count_27_io_out ? io_r_101_b : _GEN_11080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11082 = 9'h66 == r_count_27_io_out ? io_r_102_b : _GEN_11081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11083 = 9'h67 == r_count_27_io_out ? io_r_103_b : _GEN_11082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11084 = 9'h68 == r_count_27_io_out ? io_r_104_b : _GEN_11083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11085 = 9'h69 == r_count_27_io_out ? io_r_105_b : _GEN_11084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11086 = 9'h6a == r_count_27_io_out ? io_r_106_b : _GEN_11085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11087 = 9'h6b == r_count_27_io_out ? io_r_107_b : _GEN_11086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11088 = 9'h6c == r_count_27_io_out ? io_r_108_b : _GEN_11087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11089 = 9'h6d == r_count_27_io_out ? io_r_109_b : _GEN_11088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11090 = 9'h6e == r_count_27_io_out ? io_r_110_b : _GEN_11089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11091 = 9'h6f == r_count_27_io_out ? io_r_111_b : _GEN_11090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11092 = 9'h70 == r_count_27_io_out ? io_r_112_b : _GEN_11091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11093 = 9'h71 == r_count_27_io_out ? io_r_113_b : _GEN_11092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11094 = 9'h72 == r_count_27_io_out ? io_r_114_b : _GEN_11093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11095 = 9'h73 == r_count_27_io_out ? io_r_115_b : _GEN_11094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11096 = 9'h74 == r_count_27_io_out ? io_r_116_b : _GEN_11095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11097 = 9'h75 == r_count_27_io_out ? io_r_117_b : _GEN_11096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11098 = 9'h76 == r_count_27_io_out ? io_r_118_b : _GEN_11097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11099 = 9'h77 == r_count_27_io_out ? io_r_119_b : _GEN_11098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11100 = 9'h78 == r_count_27_io_out ? io_r_120_b : _GEN_11099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11101 = 9'h79 == r_count_27_io_out ? io_r_121_b : _GEN_11100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11102 = 9'h7a == r_count_27_io_out ? io_r_122_b : _GEN_11101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11103 = 9'h7b == r_count_27_io_out ? io_r_123_b : _GEN_11102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11104 = 9'h7c == r_count_27_io_out ? io_r_124_b : _GEN_11103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11105 = 9'h7d == r_count_27_io_out ? io_r_125_b : _GEN_11104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11106 = 9'h7e == r_count_27_io_out ? io_r_126_b : _GEN_11105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11107 = 9'h7f == r_count_27_io_out ? io_r_127_b : _GEN_11106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11108 = 9'h80 == r_count_27_io_out ? io_r_128_b : _GEN_11107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11109 = 9'h81 == r_count_27_io_out ? io_r_129_b : _GEN_11108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11110 = 9'h82 == r_count_27_io_out ? io_r_130_b : _GEN_11109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11111 = 9'h83 == r_count_27_io_out ? io_r_131_b : _GEN_11110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11112 = 9'h84 == r_count_27_io_out ? io_r_132_b : _GEN_11111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11113 = 9'h85 == r_count_27_io_out ? io_r_133_b : _GEN_11112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11114 = 9'h86 == r_count_27_io_out ? io_r_134_b : _GEN_11113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11115 = 9'h87 == r_count_27_io_out ? io_r_135_b : _GEN_11114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11116 = 9'h88 == r_count_27_io_out ? io_r_136_b : _GEN_11115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11117 = 9'h89 == r_count_27_io_out ? io_r_137_b : _GEN_11116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11118 = 9'h8a == r_count_27_io_out ? io_r_138_b : _GEN_11117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11119 = 9'h8b == r_count_27_io_out ? io_r_139_b : _GEN_11118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11120 = 9'h8c == r_count_27_io_out ? io_r_140_b : _GEN_11119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11121 = 9'h8d == r_count_27_io_out ? io_r_141_b : _GEN_11120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11122 = 9'h8e == r_count_27_io_out ? io_r_142_b : _GEN_11121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11123 = 9'h8f == r_count_27_io_out ? io_r_143_b : _GEN_11122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11124 = 9'h90 == r_count_27_io_out ? io_r_144_b : _GEN_11123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11125 = 9'h91 == r_count_27_io_out ? io_r_145_b : _GEN_11124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11126 = 9'h92 == r_count_27_io_out ? io_r_146_b : _GEN_11125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11127 = 9'h93 == r_count_27_io_out ? io_r_147_b : _GEN_11126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11128 = 9'h94 == r_count_27_io_out ? io_r_148_b : _GEN_11127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11129 = 9'h95 == r_count_27_io_out ? io_r_149_b : _GEN_11128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11130 = 9'h96 == r_count_27_io_out ? io_r_150_b : _GEN_11129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11131 = 9'h97 == r_count_27_io_out ? io_r_151_b : _GEN_11130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11132 = 9'h98 == r_count_27_io_out ? io_r_152_b : _GEN_11131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11133 = 9'h99 == r_count_27_io_out ? io_r_153_b : _GEN_11132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11134 = 9'h9a == r_count_27_io_out ? io_r_154_b : _GEN_11133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11135 = 9'h9b == r_count_27_io_out ? io_r_155_b : _GEN_11134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11136 = 9'h9c == r_count_27_io_out ? io_r_156_b : _GEN_11135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11137 = 9'h9d == r_count_27_io_out ? io_r_157_b : _GEN_11136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11138 = 9'h9e == r_count_27_io_out ? io_r_158_b : _GEN_11137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11139 = 9'h9f == r_count_27_io_out ? io_r_159_b : _GEN_11138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11140 = 9'ha0 == r_count_27_io_out ? io_r_160_b : _GEN_11139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11141 = 9'ha1 == r_count_27_io_out ? io_r_161_b : _GEN_11140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11142 = 9'ha2 == r_count_27_io_out ? io_r_162_b : _GEN_11141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11143 = 9'ha3 == r_count_27_io_out ? io_r_163_b : _GEN_11142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11144 = 9'ha4 == r_count_27_io_out ? io_r_164_b : _GEN_11143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11145 = 9'ha5 == r_count_27_io_out ? io_r_165_b : _GEN_11144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11146 = 9'ha6 == r_count_27_io_out ? io_r_166_b : _GEN_11145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11147 = 9'ha7 == r_count_27_io_out ? io_r_167_b : _GEN_11146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11148 = 9'ha8 == r_count_27_io_out ? io_r_168_b : _GEN_11147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11149 = 9'ha9 == r_count_27_io_out ? io_r_169_b : _GEN_11148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11150 = 9'haa == r_count_27_io_out ? io_r_170_b : _GEN_11149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11151 = 9'hab == r_count_27_io_out ? io_r_171_b : _GEN_11150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11152 = 9'hac == r_count_27_io_out ? io_r_172_b : _GEN_11151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11153 = 9'had == r_count_27_io_out ? io_r_173_b : _GEN_11152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11154 = 9'hae == r_count_27_io_out ? io_r_174_b : _GEN_11153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11155 = 9'haf == r_count_27_io_out ? io_r_175_b : _GEN_11154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11156 = 9'hb0 == r_count_27_io_out ? io_r_176_b : _GEN_11155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11157 = 9'hb1 == r_count_27_io_out ? io_r_177_b : _GEN_11156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11158 = 9'hb2 == r_count_27_io_out ? io_r_178_b : _GEN_11157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11159 = 9'hb3 == r_count_27_io_out ? io_r_179_b : _GEN_11158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11160 = 9'hb4 == r_count_27_io_out ? io_r_180_b : _GEN_11159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11161 = 9'hb5 == r_count_27_io_out ? io_r_181_b : _GEN_11160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11162 = 9'hb6 == r_count_27_io_out ? io_r_182_b : _GEN_11161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11163 = 9'hb7 == r_count_27_io_out ? io_r_183_b : _GEN_11162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11164 = 9'hb8 == r_count_27_io_out ? io_r_184_b : _GEN_11163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11165 = 9'hb9 == r_count_27_io_out ? io_r_185_b : _GEN_11164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11166 = 9'hba == r_count_27_io_out ? io_r_186_b : _GEN_11165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11167 = 9'hbb == r_count_27_io_out ? io_r_187_b : _GEN_11166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11168 = 9'hbc == r_count_27_io_out ? io_r_188_b : _GEN_11167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11169 = 9'hbd == r_count_27_io_out ? io_r_189_b : _GEN_11168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11170 = 9'hbe == r_count_27_io_out ? io_r_190_b : _GEN_11169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11171 = 9'hbf == r_count_27_io_out ? io_r_191_b : _GEN_11170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11172 = 9'hc0 == r_count_27_io_out ? io_r_192_b : _GEN_11171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11173 = 9'hc1 == r_count_27_io_out ? io_r_193_b : _GEN_11172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11174 = 9'hc2 == r_count_27_io_out ? io_r_194_b : _GEN_11173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11175 = 9'hc3 == r_count_27_io_out ? io_r_195_b : _GEN_11174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11176 = 9'hc4 == r_count_27_io_out ? io_r_196_b : _GEN_11175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11177 = 9'hc5 == r_count_27_io_out ? io_r_197_b : _GEN_11176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11178 = 9'hc6 == r_count_27_io_out ? io_r_198_b : _GEN_11177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11179 = 9'hc7 == r_count_27_io_out ? io_r_199_b : _GEN_11178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11180 = 9'hc8 == r_count_27_io_out ? io_r_200_b : _GEN_11179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11181 = 9'hc9 == r_count_27_io_out ? io_r_201_b : _GEN_11180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11182 = 9'hca == r_count_27_io_out ? io_r_202_b : _GEN_11181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11183 = 9'hcb == r_count_27_io_out ? io_r_203_b : _GEN_11182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11184 = 9'hcc == r_count_27_io_out ? io_r_204_b : _GEN_11183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11185 = 9'hcd == r_count_27_io_out ? io_r_205_b : _GEN_11184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11186 = 9'hce == r_count_27_io_out ? io_r_206_b : _GEN_11185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11187 = 9'hcf == r_count_27_io_out ? io_r_207_b : _GEN_11186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11188 = 9'hd0 == r_count_27_io_out ? io_r_208_b : _GEN_11187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11189 = 9'hd1 == r_count_27_io_out ? io_r_209_b : _GEN_11188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11190 = 9'hd2 == r_count_27_io_out ? io_r_210_b : _GEN_11189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11191 = 9'hd3 == r_count_27_io_out ? io_r_211_b : _GEN_11190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11192 = 9'hd4 == r_count_27_io_out ? io_r_212_b : _GEN_11191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11193 = 9'hd5 == r_count_27_io_out ? io_r_213_b : _GEN_11192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11194 = 9'hd6 == r_count_27_io_out ? io_r_214_b : _GEN_11193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11195 = 9'hd7 == r_count_27_io_out ? io_r_215_b : _GEN_11194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11196 = 9'hd8 == r_count_27_io_out ? io_r_216_b : _GEN_11195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11197 = 9'hd9 == r_count_27_io_out ? io_r_217_b : _GEN_11196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11198 = 9'hda == r_count_27_io_out ? io_r_218_b : _GEN_11197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11199 = 9'hdb == r_count_27_io_out ? io_r_219_b : _GEN_11198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11200 = 9'hdc == r_count_27_io_out ? io_r_220_b : _GEN_11199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11201 = 9'hdd == r_count_27_io_out ? io_r_221_b : _GEN_11200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11202 = 9'hde == r_count_27_io_out ? io_r_222_b : _GEN_11201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11203 = 9'hdf == r_count_27_io_out ? io_r_223_b : _GEN_11202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11204 = 9'he0 == r_count_27_io_out ? io_r_224_b : _GEN_11203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11205 = 9'he1 == r_count_27_io_out ? io_r_225_b : _GEN_11204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11206 = 9'he2 == r_count_27_io_out ? io_r_226_b : _GEN_11205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11207 = 9'he3 == r_count_27_io_out ? io_r_227_b : _GEN_11206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11208 = 9'he4 == r_count_27_io_out ? io_r_228_b : _GEN_11207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11209 = 9'he5 == r_count_27_io_out ? io_r_229_b : _GEN_11208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11210 = 9'he6 == r_count_27_io_out ? io_r_230_b : _GEN_11209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11211 = 9'he7 == r_count_27_io_out ? io_r_231_b : _GEN_11210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11212 = 9'he8 == r_count_27_io_out ? io_r_232_b : _GEN_11211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11213 = 9'he9 == r_count_27_io_out ? io_r_233_b : _GEN_11212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11214 = 9'hea == r_count_27_io_out ? io_r_234_b : _GEN_11213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11215 = 9'heb == r_count_27_io_out ? io_r_235_b : _GEN_11214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11216 = 9'hec == r_count_27_io_out ? io_r_236_b : _GEN_11215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11217 = 9'hed == r_count_27_io_out ? io_r_237_b : _GEN_11216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11218 = 9'hee == r_count_27_io_out ? io_r_238_b : _GEN_11217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11219 = 9'hef == r_count_27_io_out ? io_r_239_b : _GEN_11218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11220 = 9'hf0 == r_count_27_io_out ? io_r_240_b : _GEN_11219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11221 = 9'hf1 == r_count_27_io_out ? io_r_241_b : _GEN_11220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11222 = 9'hf2 == r_count_27_io_out ? io_r_242_b : _GEN_11221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11223 = 9'hf3 == r_count_27_io_out ? io_r_243_b : _GEN_11222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11224 = 9'hf4 == r_count_27_io_out ? io_r_244_b : _GEN_11223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11225 = 9'hf5 == r_count_27_io_out ? io_r_245_b : _GEN_11224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11226 = 9'hf6 == r_count_27_io_out ? io_r_246_b : _GEN_11225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11227 = 9'hf7 == r_count_27_io_out ? io_r_247_b : _GEN_11226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11228 = 9'hf8 == r_count_27_io_out ? io_r_248_b : _GEN_11227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11229 = 9'hf9 == r_count_27_io_out ? io_r_249_b : _GEN_11228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11230 = 9'hfa == r_count_27_io_out ? io_r_250_b : _GEN_11229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11231 = 9'hfb == r_count_27_io_out ? io_r_251_b : _GEN_11230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11232 = 9'hfc == r_count_27_io_out ? io_r_252_b : _GEN_11231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11233 = 9'hfd == r_count_27_io_out ? io_r_253_b : _GEN_11232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11234 = 9'hfe == r_count_27_io_out ? io_r_254_b : _GEN_11233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11235 = 9'hff == r_count_27_io_out ? io_r_255_b : _GEN_11234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11236 = 9'h100 == r_count_27_io_out ? io_r_256_b : _GEN_11235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11237 = 9'h101 == r_count_27_io_out ? io_r_257_b : _GEN_11236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11238 = 9'h102 == r_count_27_io_out ? io_r_258_b : _GEN_11237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11239 = 9'h103 == r_count_27_io_out ? io_r_259_b : _GEN_11238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11240 = 9'h104 == r_count_27_io_out ? io_r_260_b : _GEN_11239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11241 = 9'h105 == r_count_27_io_out ? io_r_261_b : _GEN_11240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11242 = 9'h106 == r_count_27_io_out ? io_r_262_b : _GEN_11241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11243 = 9'h107 == r_count_27_io_out ? io_r_263_b : _GEN_11242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11244 = 9'h108 == r_count_27_io_out ? io_r_264_b : _GEN_11243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11245 = 9'h109 == r_count_27_io_out ? io_r_265_b : _GEN_11244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11246 = 9'h10a == r_count_27_io_out ? io_r_266_b : _GEN_11245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11247 = 9'h10b == r_count_27_io_out ? io_r_267_b : _GEN_11246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11248 = 9'h10c == r_count_27_io_out ? io_r_268_b : _GEN_11247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11249 = 9'h10d == r_count_27_io_out ? io_r_269_b : _GEN_11248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11250 = 9'h10e == r_count_27_io_out ? io_r_270_b : _GEN_11249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11251 = 9'h10f == r_count_27_io_out ? io_r_271_b : _GEN_11250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11252 = 9'h110 == r_count_27_io_out ? io_r_272_b : _GEN_11251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11253 = 9'h111 == r_count_27_io_out ? io_r_273_b : _GEN_11252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11254 = 9'h112 == r_count_27_io_out ? io_r_274_b : _GEN_11253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11255 = 9'h113 == r_count_27_io_out ? io_r_275_b : _GEN_11254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11256 = 9'h114 == r_count_27_io_out ? io_r_276_b : _GEN_11255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11257 = 9'h115 == r_count_27_io_out ? io_r_277_b : _GEN_11256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11258 = 9'h116 == r_count_27_io_out ? io_r_278_b : _GEN_11257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11259 = 9'h117 == r_count_27_io_out ? io_r_279_b : _GEN_11258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11260 = 9'h118 == r_count_27_io_out ? io_r_280_b : _GEN_11259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11261 = 9'h119 == r_count_27_io_out ? io_r_281_b : _GEN_11260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11262 = 9'h11a == r_count_27_io_out ? io_r_282_b : _GEN_11261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11263 = 9'h11b == r_count_27_io_out ? io_r_283_b : _GEN_11262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11264 = 9'h11c == r_count_27_io_out ? io_r_284_b : _GEN_11263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11265 = 9'h11d == r_count_27_io_out ? io_r_285_b : _GEN_11264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11266 = 9'h11e == r_count_27_io_out ? io_r_286_b : _GEN_11265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11267 = 9'h11f == r_count_27_io_out ? io_r_287_b : _GEN_11266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11268 = 9'h120 == r_count_27_io_out ? io_r_288_b : _GEN_11267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11269 = 9'h121 == r_count_27_io_out ? io_r_289_b : _GEN_11268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11270 = 9'h122 == r_count_27_io_out ? io_r_290_b : _GEN_11269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11271 = 9'h123 == r_count_27_io_out ? io_r_291_b : _GEN_11270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11272 = 9'h124 == r_count_27_io_out ? io_r_292_b : _GEN_11271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11273 = 9'h125 == r_count_27_io_out ? io_r_293_b : _GEN_11272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11274 = 9'h126 == r_count_27_io_out ? io_r_294_b : _GEN_11273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11275 = 9'h127 == r_count_27_io_out ? io_r_295_b : _GEN_11274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11276 = 9'h128 == r_count_27_io_out ? io_r_296_b : _GEN_11275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11277 = 9'h129 == r_count_27_io_out ? io_r_297_b : _GEN_11276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11278 = 9'h12a == r_count_27_io_out ? io_r_298_b : _GEN_11277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11279 = 9'h12b == r_count_27_io_out ? io_r_299_b : _GEN_11278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11280 = 9'h12c == r_count_27_io_out ? io_r_300_b : _GEN_11279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11281 = 9'h12d == r_count_27_io_out ? io_r_301_b : _GEN_11280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11282 = 9'h12e == r_count_27_io_out ? io_r_302_b : _GEN_11281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11283 = 9'h12f == r_count_27_io_out ? io_r_303_b : _GEN_11282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11284 = 9'h130 == r_count_27_io_out ? io_r_304_b : _GEN_11283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11285 = 9'h131 == r_count_27_io_out ? io_r_305_b : _GEN_11284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11286 = 9'h132 == r_count_27_io_out ? io_r_306_b : _GEN_11285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11287 = 9'h133 == r_count_27_io_out ? io_r_307_b : _GEN_11286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11288 = 9'h134 == r_count_27_io_out ? io_r_308_b : _GEN_11287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11289 = 9'h135 == r_count_27_io_out ? io_r_309_b : _GEN_11288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11290 = 9'h136 == r_count_27_io_out ? io_r_310_b : _GEN_11289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11291 = 9'h137 == r_count_27_io_out ? io_r_311_b : _GEN_11290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11292 = 9'h138 == r_count_27_io_out ? io_r_312_b : _GEN_11291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11293 = 9'h139 == r_count_27_io_out ? io_r_313_b : _GEN_11292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11294 = 9'h13a == r_count_27_io_out ? io_r_314_b : _GEN_11293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11295 = 9'h13b == r_count_27_io_out ? io_r_315_b : _GEN_11294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11296 = 9'h13c == r_count_27_io_out ? io_r_316_b : _GEN_11295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11297 = 9'h13d == r_count_27_io_out ? io_r_317_b : _GEN_11296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11298 = 9'h13e == r_count_27_io_out ? io_r_318_b : _GEN_11297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11299 = 9'h13f == r_count_27_io_out ? io_r_319_b : _GEN_11298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11300 = 9'h140 == r_count_27_io_out ? io_r_320_b : _GEN_11299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11301 = 9'h141 == r_count_27_io_out ? io_r_321_b : _GEN_11300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11302 = 9'h142 == r_count_27_io_out ? io_r_322_b : _GEN_11301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11303 = 9'h143 == r_count_27_io_out ? io_r_323_b : _GEN_11302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11304 = 9'h144 == r_count_27_io_out ? io_r_324_b : _GEN_11303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11305 = 9'h145 == r_count_27_io_out ? io_r_325_b : _GEN_11304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11306 = 9'h146 == r_count_27_io_out ? io_r_326_b : _GEN_11305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11307 = 9'h147 == r_count_27_io_out ? io_r_327_b : _GEN_11306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11308 = 9'h148 == r_count_27_io_out ? io_r_328_b : _GEN_11307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11309 = 9'h149 == r_count_27_io_out ? io_r_329_b : _GEN_11308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11310 = 9'h14a == r_count_27_io_out ? io_r_330_b : _GEN_11309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11311 = 9'h14b == r_count_27_io_out ? io_r_331_b : _GEN_11310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11312 = 9'h14c == r_count_27_io_out ? io_r_332_b : _GEN_11311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11313 = 9'h14d == r_count_27_io_out ? io_r_333_b : _GEN_11312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11314 = 9'h14e == r_count_27_io_out ? io_r_334_b : _GEN_11313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11315 = 9'h14f == r_count_27_io_out ? io_r_335_b : _GEN_11314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11316 = 9'h150 == r_count_27_io_out ? io_r_336_b : _GEN_11315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11317 = 9'h151 == r_count_27_io_out ? io_r_337_b : _GEN_11316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11318 = 9'h152 == r_count_27_io_out ? io_r_338_b : _GEN_11317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11319 = 9'h153 == r_count_27_io_out ? io_r_339_b : _GEN_11318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11320 = 9'h154 == r_count_27_io_out ? io_r_340_b : _GEN_11319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11321 = 9'h155 == r_count_27_io_out ? io_r_341_b : _GEN_11320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11322 = 9'h156 == r_count_27_io_out ? io_r_342_b : _GEN_11321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11323 = 9'h157 == r_count_27_io_out ? io_r_343_b : _GEN_11322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11324 = 9'h158 == r_count_27_io_out ? io_r_344_b : _GEN_11323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11325 = 9'h159 == r_count_27_io_out ? io_r_345_b : _GEN_11324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11326 = 9'h15a == r_count_27_io_out ? io_r_346_b : _GEN_11325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11327 = 9'h15b == r_count_27_io_out ? io_r_347_b : _GEN_11326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11328 = 9'h15c == r_count_27_io_out ? io_r_348_b : _GEN_11327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11329 = 9'h15d == r_count_27_io_out ? io_r_349_b : _GEN_11328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11330 = 9'h15e == r_count_27_io_out ? io_r_350_b : _GEN_11329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11331 = 9'h15f == r_count_27_io_out ? io_r_351_b : _GEN_11330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11332 = 9'h160 == r_count_27_io_out ? io_r_352_b : _GEN_11331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11333 = 9'h161 == r_count_27_io_out ? io_r_353_b : _GEN_11332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11334 = 9'h162 == r_count_27_io_out ? io_r_354_b : _GEN_11333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11335 = 9'h163 == r_count_27_io_out ? io_r_355_b : _GEN_11334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11336 = 9'h164 == r_count_27_io_out ? io_r_356_b : _GEN_11335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11337 = 9'h165 == r_count_27_io_out ? io_r_357_b : _GEN_11336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11338 = 9'h166 == r_count_27_io_out ? io_r_358_b : _GEN_11337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11339 = 9'h167 == r_count_27_io_out ? io_r_359_b : _GEN_11338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11340 = 9'h168 == r_count_27_io_out ? io_r_360_b : _GEN_11339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11341 = 9'h169 == r_count_27_io_out ? io_r_361_b : _GEN_11340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11342 = 9'h16a == r_count_27_io_out ? io_r_362_b : _GEN_11341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11343 = 9'h16b == r_count_27_io_out ? io_r_363_b : _GEN_11342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11344 = 9'h16c == r_count_27_io_out ? io_r_364_b : _GEN_11343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11345 = 9'h16d == r_count_27_io_out ? io_r_365_b : _GEN_11344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11346 = 9'h16e == r_count_27_io_out ? io_r_366_b : _GEN_11345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11347 = 9'h16f == r_count_27_io_out ? io_r_367_b : _GEN_11346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11348 = 9'h170 == r_count_27_io_out ? io_r_368_b : _GEN_11347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11349 = 9'h171 == r_count_27_io_out ? io_r_369_b : _GEN_11348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11350 = 9'h172 == r_count_27_io_out ? io_r_370_b : _GEN_11349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11351 = 9'h173 == r_count_27_io_out ? io_r_371_b : _GEN_11350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11352 = 9'h174 == r_count_27_io_out ? io_r_372_b : _GEN_11351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11353 = 9'h175 == r_count_27_io_out ? io_r_373_b : _GEN_11352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11354 = 9'h176 == r_count_27_io_out ? io_r_374_b : _GEN_11353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11355 = 9'h177 == r_count_27_io_out ? io_r_375_b : _GEN_11354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11356 = 9'h178 == r_count_27_io_out ? io_r_376_b : _GEN_11355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11357 = 9'h179 == r_count_27_io_out ? io_r_377_b : _GEN_11356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11358 = 9'h17a == r_count_27_io_out ? io_r_378_b : _GEN_11357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11359 = 9'h17b == r_count_27_io_out ? io_r_379_b : _GEN_11358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11360 = 9'h17c == r_count_27_io_out ? io_r_380_b : _GEN_11359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11361 = 9'h17d == r_count_27_io_out ? io_r_381_b : _GEN_11360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11362 = 9'h17e == r_count_27_io_out ? io_r_382_b : _GEN_11361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11363 = 9'h17f == r_count_27_io_out ? io_r_383_b : _GEN_11362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11364 = 9'h180 == r_count_27_io_out ? io_r_384_b : _GEN_11363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11365 = 9'h181 == r_count_27_io_out ? io_r_385_b : _GEN_11364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11366 = 9'h182 == r_count_27_io_out ? io_r_386_b : _GEN_11365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11367 = 9'h183 == r_count_27_io_out ? io_r_387_b : _GEN_11366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11368 = 9'h184 == r_count_27_io_out ? io_r_388_b : _GEN_11367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11369 = 9'h185 == r_count_27_io_out ? io_r_389_b : _GEN_11368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11370 = 9'h186 == r_count_27_io_out ? io_r_390_b : _GEN_11369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11371 = 9'h187 == r_count_27_io_out ? io_r_391_b : _GEN_11370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11372 = 9'h188 == r_count_27_io_out ? io_r_392_b : _GEN_11371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11373 = 9'h189 == r_count_27_io_out ? io_r_393_b : _GEN_11372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11374 = 9'h18a == r_count_27_io_out ? io_r_394_b : _GEN_11373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11375 = 9'h18b == r_count_27_io_out ? io_r_395_b : _GEN_11374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11376 = 9'h18c == r_count_27_io_out ? io_r_396_b : _GEN_11375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11377 = 9'h18d == r_count_27_io_out ? io_r_397_b : _GEN_11376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11378 = 9'h18e == r_count_27_io_out ? io_r_398_b : _GEN_11377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11381 = 9'h1 == r_count_28_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11382 = 9'h2 == r_count_28_io_out ? io_r_2_b : _GEN_11381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11383 = 9'h3 == r_count_28_io_out ? io_r_3_b : _GEN_11382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11384 = 9'h4 == r_count_28_io_out ? io_r_4_b : _GEN_11383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11385 = 9'h5 == r_count_28_io_out ? io_r_5_b : _GEN_11384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11386 = 9'h6 == r_count_28_io_out ? io_r_6_b : _GEN_11385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11387 = 9'h7 == r_count_28_io_out ? io_r_7_b : _GEN_11386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11388 = 9'h8 == r_count_28_io_out ? io_r_8_b : _GEN_11387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11389 = 9'h9 == r_count_28_io_out ? io_r_9_b : _GEN_11388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11390 = 9'ha == r_count_28_io_out ? io_r_10_b : _GEN_11389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11391 = 9'hb == r_count_28_io_out ? io_r_11_b : _GEN_11390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11392 = 9'hc == r_count_28_io_out ? io_r_12_b : _GEN_11391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11393 = 9'hd == r_count_28_io_out ? io_r_13_b : _GEN_11392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11394 = 9'he == r_count_28_io_out ? io_r_14_b : _GEN_11393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11395 = 9'hf == r_count_28_io_out ? io_r_15_b : _GEN_11394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11396 = 9'h10 == r_count_28_io_out ? io_r_16_b : _GEN_11395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11397 = 9'h11 == r_count_28_io_out ? io_r_17_b : _GEN_11396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11398 = 9'h12 == r_count_28_io_out ? io_r_18_b : _GEN_11397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11399 = 9'h13 == r_count_28_io_out ? io_r_19_b : _GEN_11398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11400 = 9'h14 == r_count_28_io_out ? io_r_20_b : _GEN_11399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11401 = 9'h15 == r_count_28_io_out ? io_r_21_b : _GEN_11400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11402 = 9'h16 == r_count_28_io_out ? io_r_22_b : _GEN_11401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11403 = 9'h17 == r_count_28_io_out ? io_r_23_b : _GEN_11402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11404 = 9'h18 == r_count_28_io_out ? io_r_24_b : _GEN_11403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11405 = 9'h19 == r_count_28_io_out ? io_r_25_b : _GEN_11404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11406 = 9'h1a == r_count_28_io_out ? io_r_26_b : _GEN_11405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11407 = 9'h1b == r_count_28_io_out ? io_r_27_b : _GEN_11406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11408 = 9'h1c == r_count_28_io_out ? io_r_28_b : _GEN_11407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11409 = 9'h1d == r_count_28_io_out ? io_r_29_b : _GEN_11408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11410 = 9'h1e == r_count_28_io_out ? io_r_30_b : _GEN_11409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11411 = 9'h1f == r_count_28_io_out ? io_r_31_b : _GEN_11410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11412 = 9'h20 == r_count_28_io_out ? io_r_32_b : _GEN_11411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11413 = 9'h21 == r_count_28_io_out ? io_r_33_b : _GEN_11412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11414 = 9'h22 == r_count_28_io_out ? io_r_34_b : _GEN_11413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11415 = 9'h23 == r_count_28_io_out ? io_r_35_b : _GEN_11414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11416 = 9'h24 == r_count_28_io_out ? io_r_36_b : _GEN_11415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11417 = 9'h25 == r_count_28_io_out ? io_r_37_b : _GEN_11416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11418 = 9'h26 == r_count_28_io_out ? io_r_38_b : _GEN_11417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11419 = 9'h27 == r_count_28_io_out ? io_r_39_b : _GEN_11418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11420 = 9'h28 == r_count_28_io_out ? io_r_40_b : _GEN_11419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11421 = 9'h29 == r_count_28_io_out ? io_r_41_b : _GEN_11420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11422 = 9'h2a == r_count_28_io_out ? io_r_42_b : _GEN_11421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11423 = 9'h2b == r_count_28_io_out ? io_r_43_b : _GEN_11422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11424 = 9'h2c == r_count_28_io_out ? io_r_44_b : _GEN_11423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11425 = 9'h2d == r_count_28_io_out ? io_r_45_b : _GEN_11424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11426 = 9'h2e == r_count_28_io_out ? io_r_46_b : _GEN_11425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11427 = 9'h2f == r_count_28_io_out ? io_r_47_b : _GEN_11426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11428 = 9'h30 == r_count_28_io_out ? io_r_48_b : _GEN_11427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11429 = 9'h31 == r_count_28_io_out ? io_r_49_b : _GEN_11428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11430 = 9'h32 == r_count_28_io_out ? io_r_50_b : _GEN_11429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11431 = 9'h33 == r_count_28_io_out ? io_r_51_b : _GEN_11430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11432 = 9'h34 == r_count_28_io_out ? io_r_52_b : _GEN_11431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11433 = 9'h35 == r_count_28_io_out ? io_r_53_b : _GEN_11432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11434 = 9'h36 == r_count_28_io_out ? io_r_54_b : _GEN_11433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11435 = 9'h37 == r_count_28_io_out ? io_r_55_b : _GEN_11434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11436 = 9'h38 == r_count_28_io_out ? io_r_56_b : _GEN_11435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11437 = 9'h39 == r_count_28_io_out ? io_r_57_b : _GEN_11436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11438 = 9'h3a == r_count_28_io_out ? io_r_58_b : _GEN_11437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11439 = 9'h3b == r_count_28_io_out ? io_r_59_b : _GEN_11438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11440 = 9'h3c == r_count_28_io_out ? io_r_60_b : _GEN_11439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11441 = 9'h3d == r_count_28_io_out ? io_r_61_b : _GEN_11440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11442 = 9'h3e == r_count_28_io_out ? io_r_62_b : _GEN_11441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11443 = 9'h3f == r_count_28_io_out ? io_r_63_b : _GEN_11442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11444 = 9'h40 == r_count_28_io_out ? io_r_64_b : _GEN_11443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11445 = 9'h41 == r_count_28_io_out ? io_r_65_b : _GEN_11444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11446 = 9'h42 == r_count_28_io_out ? io_r_66_b : _GEN_11445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11447 = 9'h43 == r_count_28_io_out ? io_r_67_b : _GEN_11446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11448 = 9'h44 == r_count_28_io_out ? io_r_68_b : _GEN_11447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11449 = 9'h45 == r_count_28_io_out ? io_r_69_b : _GEN_11448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11450 = 9'h46 == r_count_28_io_out ? io_r_70_b : _GEN_11449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11451 = 9'h47 == r_count_28_io_out ? io_r_71_b : _GEN_11450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11452 = 9'h48 == r_count_28_io_out ? io_r_72_b : _GEN_11451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11453 = 9'h49 == r_count_28_io_out ? io_r_73_b : _GEN_11452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11454 = 9'h4a == r_count_28_io_out ? io_r_74_b : _GEN_11453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11455 = 9'h4b == r_count_28_io_out ? io_r_75_b : _GEN_11454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11456 = 9'h4c == r_count_28_io_out ? io_r_76_b : _GEN_11455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11457 = 9'h4d == r_count_28_io_out ? io_r_77_b : _GEN_11456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11458 = 9'h4e == r_count_28_io_out ? io_r_78_b : _GEN_11457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11459 = 9'h4f == r_count_28_io_out ? io_r_79_b : _GEN_11458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11460 = 9'h50 == r_count_28_io_out ? io_r_80_b : _GEN_11459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11461 = 9'h51 == r_count_28_io_out ? io_r_81_b : _GEN_11460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11462 = 9'h52 == r_count_28_io_out ? io_r_82_b : _GEN_11461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11463 = 9'h53 == r_count_28_io_out ? io_r_83_b : _GEN_11462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11464 = 9'h54 == r_count_28_io_out ? io_r_84_b : _GEN_11463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11465 = 9'h55 == r_count_28_io_out ? io_r_85_b : _GEN_11464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11466 = 9'h56 == r_count_28_io_out ? io_r_86_b : _GEN_11465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11467 = 9'h57 == r_count_28_io_out ? io_r_87_b : _GEN_11466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11468 = 9'h58 == r_count_28_io_out ? io_r_88_b : _GEN_11467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11469 = 9'h59 == r_count_28_io_out ? io_r_89_b : _GEN_11468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11470 = 9'h5a == r_count_28_io_out ? io_r_90_b : _GEN_11469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11471 = 9'h5b == r_count_28_io_out ? io_r_91_b : _GEN_11470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11472 = 9'h5c == r_count_28_io_out ? io_r_92_b : _GEN_11471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11473 = 9'h5d == r_count_28_io_out ? io_r_93_b : _GEN_11472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11474 = 9'h5e == r_count_28_io_out ? io_r_94_b : _GEN_11473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11475 = 9'h5f == r_count_28_io_out ? io_r_95_b : _GEN_11474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11476 = 9'h60 == r_count_28_io_out ? io_r_96_b : _GEN_11475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11477 = 9'h61 == r_count_28_io_out ? io_r_97_b : _GEN_11476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11478 = 9'h62 == r_count_28_io_out ? io_r_98_b : _GEN_11477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11479 = 9'h63 == r_count_28_io_out ? io_r_99_b : _GEN_11478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11480 = 9'h64 == r_count_28_io_out ? io_r_100_b : _GEN_11479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11481 = 9'h65 == r_count_28_io_out ? io_r_101_b : _GEN_11480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11482 = 9'h66 == r_count_28_io_out ? io_r_102_b : _GEN_11481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11483 = 9'h67 == r_count_28_io_out ? io_r_103_b : _GEN_11482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11484 = 9'h68 == r_count_28_io_out ? io_r_104_b : _GEN_11483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11485 = 9'h69 == r_count_28_io_out ? io_r_105_b : _GEN_11484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11486 = 9'h6a == r_count_28_io_out ? io_r_106_b : _GEN_11485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11487 = 9'h6b == r_count_28_io_out ? io_r_107_b : _GEN_11486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11488 = 9'h6c == r_count_28_io_out ? io_r_108_b : _GEN_11487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11489 = 9'h6d == r_count_28_io_out ? io_r_109_b : _GEN_11488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11490 = 9'h6e == r_count_28_io_out ? io_r_110_b : _GEN_11489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11491 = 9'h6f == r_count_28_io_out ? io_r_111_b : _GEN_11490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11492 = 9'h70 == r_count_28_io_out ? io_r_112_b : _GEN_11491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11493 = 9'h71 == r_count_28_io_out ? io_r_113_b : _GEN_11492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11494 = 9'h72 == r_count_28_io_out ? io_r_114_b : _GEN_11493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11495 = 9'h73 == r_count_28_io_out ? io_r_115_b : _GEN_11494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11496 = 9'h74 == r_count_28_io_out ? io_r_116_b : _GEN_11495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11497 = 9'h75 == r_count_28_io_out ? io_r_117_b : _GEN_11496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11498 = 9'h76 == r_count_28_io_out ? io_r_118_b : _GEN_11497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11499 = 9'h77 == r_count_28_io_out ? io_r_119_b : _GEN_11498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11500 = 9'h78 == r_count_28_io_out ? io_r_120_b : _GEN_11499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11501 = 9'h79 == r_count_28_io_out ? io_r_121_b : _GEN_11500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11502 = 9'h7a == r_count_28_io_out ? io_r_122_b : _GEN_11501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11503 = 9'h7b == r_count_28_io_out ? io_r_123_b : _GEN_11502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11504 = 9'h7c == r_count_28_io_out ? io_r_124_b : _GEN_11503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11505 = 9'h7d == r_count_28_io_out ? io_r_125_b : _GEN_11504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11506 = 9'h7e == r_count_28_io_out ? io_r_126_b : _GEN_11505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11507 = 9'h7f == r_count_28_io_out ? io_r_127_b : _GEN_11506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11508 = 9'h80 == r_count_28_io_out ? io_r_128_b : _GEN_11507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11509 = 9'h81 == r_count_28_io_out ? io_r_129_b : _GEN_11508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11510 = 9'h82 == r_count_28_io_out ? io_r_130_b : _GEN_11509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11511 = 9'h83 == r_count_28_io_out ? io_r_131_b : _GEN_11510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11512 = 9'h84 == r_count_28_io_out ? io_r_132_b : _GEN_11511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11513 = 9'h85 == r_count_28_io_out ? io_r_133_b : _GEN_11512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11514 = 9'h86 == r_count_28_io_out ? io_r_134_b : _GEN_11513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11515 = 9'h87 == r_count_28_io_out ? io_r_135_b : _GEN_11514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11516 = 9'h88 == r_count_28_io_out ? io_r_136_b : _GEN_11515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11517 = 9'h89 == r_count_28_io_out ? io_r_137_b : _GEN_11516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11518 = 9'h8a == r_count_28_io_out ? io_r_138_b : _GEN_11517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11519 = 9'h8b == r_count_28_io_out ? io_r_139_b : _GEN_11518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11520 = 9'h8c == r_count_28_io_out ? io_r_140_b : _GEN_11519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11521 = 9'h8d == r_count_28_io_out ? io_r_141_b : _GEN_11520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11522 = 9'h8e == r_count_28_io_out ? io_r_142_b : _GEN_11521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11523 = 9'h8f == r_count_28_io_out ? io_r_143_b : _GEN_11522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11524 = 9'h90 == r_count_28_io_out ? io_r_144_b : _GEN_11523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11525 = 9'h91 == r_count_28_io_out ? io_r_145_b : _GEN_11524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11526 = 9'h92 == r_count_28_io_out ? io_r_146_b : _GEN_11525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11527 = 9'h93 == r_count_28_io_out ? io_r_147_b : _GEN_11526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11528 = 9'h94 == r_count_28_io_out ? io_r_148_b : _GEN_11527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11529 = 9'h95 == r_count_28_io_out ? io_r_149_b : _GEN_11528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11530 = 9'h96 == r_count_28_io_out ? io_r_150_b : _GEN_11529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11531 = 9'h97 == r_count_28_io_out ? io_r_151_b : _GEN_11530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11532 = 9'h98 == r_count_28_io_out ? io_r_152_b : _GEN_11531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11533 = 9'h99 == r_count_28_io_out ? io_r_153_b : _GEN_11532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11534 = 9'h9a == r_count_28_io_out ? io_r_154_b : _GEN_11533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11535 = 9'h9b == r_count_28_io_out ? io_r_155_b : _GEN_11534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11536 = 9'h9c == r_count_28_io_out ? io_r_156_b : _GEN_11535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11537 = 9'h9d == r_count_28_io_out ? io_r_157_b : _GEN_11536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11538 = 9'h9e == r_count_28_io_out ? io_r_158_b : _GEN_11537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11539 = 9'h9f == r_count_28_io_out ? io_r_159_b : _GEN_11538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11540 = 9'ha0 == r_count_28_io_out ? io_r_160_b : _GEN_11539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11541 = 9'ha1 == r_count_28_io_out ? io_r_161_b : _GEN_11540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11542 = 9'ha2 == r_count_28_io_out ? io_r_162_b : _GEN_11541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11543 = 9'ha3 == r_count_28_io_out ? io_r_163_b : _GEN_11542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11544 = 9'ha4 == r_count_28_io_out ? io_r_164_b : _GEN_11543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11545 = 9'ha5 == r_count_28_io_out ? io_r_165_b : _GEN_11544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11546 = 9'ha6 == r_count_28_io_out ? io_r_166_b : _GEN_11545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11547 = 9'ha7 == r_count_28_io_out ? io_r_167_b : _GEN_11546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11548 = 9'ha8 == r_count_28_io_out ? io_r_168_b : _GEN_11547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11549 = 9'ha9 == r_count_28_io_out ? io_r_169_b : _GEN_11548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11550 = 9'haa == r_count_28_io_out ? io_r_170_b : _GEN_11549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11551 = 9'hab == r_count_28_io_out ? io_r_171_b : _GEN_11550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11552 = 9'hac == r_count_28_io_out ? io_r_172_b : _GEN_11551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11553 = 9'had == r_count_28_io_out ? io_r_173_b : _GEN_11552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11554 = 9'hae == r_count_28_io_out ? io_r_174_b : _GEN_11553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11555 = 9'haf == r_count_28_io_out ? io_r_175_b : _GEN_11554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11556 = 9'hb0 == r_count_28_io_out ? io_r_176_b : _GEN_11555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11557 = 9'hb1 == r_count_28_io_out ? io_r_177_b : _GEN_11556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11558 = 9'hb2 == r_count_28_io_out ? io_r_178_b : _GEN_11557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11559 = 9'hb3 == r_count_28_io_out ? io_r_179_b : _GEN_11558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11560 = 9'hb4 == r_count_28_io_out ? io_r_180_b : _GEN_11559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11561 = 9'hb5 == r_count_28_io_out ? io_r_181_b : _GEN_11560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11562 = 9'hb6 == r_count_28_io_out ? io_r_182_b : _GEN_11561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11563 = 9'hb7 == r_count_28_io_out ? io_r_183_b : _GEN_11562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11564 = 9'hb8 == r_count_28_io_out ? io_r_184_b : _GEN_11563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11565 = 9'hb9 == r_count_28_io_out ? io_r_185_b : _GEN_11564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11566 = 9'hba == r_count_28_io_out ? io_r_186_b : _GEN_11565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11567 = 9'hbb == r_count_28_io_out ? io_r_187_b : _GEN_11566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11568 = 9'hbc == r_count_28_io_out ? io_r_188_b : _GEN_11567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11569 = 9'hbd == r_count_28_io_out ? io_r_189_b : _GEN_11568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11570 = 9'hbe == r_count_28_io_out ? io_r_190_b : _GEN_11569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11571 = 9'hbf == r_count_28_io_out ? io_r_191_b : _GEN_11570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11572 = 9'hc0 == r_count_28_io_out ? io_r_192_b : _GEN_11571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11573 = 9'hc1 == r_count_28_io_out ? io_r_193_b : _GEN_11572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11574 = 9'hc2 == r_count_28_io_out ? io_r_194_b : _GEN_11573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11575 = 9'hc3 == r_count_28_io_out ? io_r_195_b : _GEN_11574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11576 = 9'hc4 == r_count_28_io_out ? io_r_196_b : _GEN_11575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11577 = 9'hc5 == r_count_28_io_out ? io_r_197_b : _GEN_11576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11578 = 9'hc6 == r_count_28_io_out ? io_r_198_b : _GEN_11577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11579 = 9'hc7 == r_count_28_io_out ? io_r_199_b : _GEN_11578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11580 = 9'hc8 == r_count_28_io_out ? io_r_200_b : _GEN_11579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11581 = 9'hc9 == r_count_28_io_out ? io_r_201_b : _GEN_11580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11582 = 9'hca == r_count_28_io_out ? io_r_202_b : _GEN_11581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11583 = 9'hcb == r_count_28_io_out ? io_r_203_b : _GEN_11582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11584 = 9'hcc == r_count_28_io_out ? io_r_204_b : _GEN_11583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11585 = 9'hcd == r_count_28_io_out ? io_r_205_b : _GEN_11584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11586 = 9'hce == r_count_28_io_out ? io_r_206_b : _GEN_11585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11587 = 9'hcf == r_count_28_io_out ? io_r_207_b : _GEN_11586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11588 = 9'hd0 == r_count_28_io_out ? io_r_208_b : _GEN_11587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11589 = 9'hd1 == r_count_28_io_out ? io_r_209_b : _GEN_11588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11590 = 9'hd2 == r_count_28_io_out ? io_r_210_b : _GEN_11589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11591 = 9'hd3 == r_count_28_io_out ? io_r_211_b : _GEN_11590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11592 = 9'hd4 == r_count_28_io_out ? io_r_212_b : _GEN_11591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11593 = 9'hd5 == r_count_28_io_out ? io_r_213_b : _GEN_11592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11594 = 9'hd6 == r_count_28_io_out ? io_r_214_b : _GEN_11593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11595 = 9'hd7 == r_count_28_io_out ? io_r_215_b : _GEN_11594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11596 = 9'hd8 == r_count_28_io_out ? io_r_216_b : _GEN_11595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11597 = 9'hd9 == r_count_28_io_out ? io_r_217_b : _GEN_11596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11598 = 9'hda == r_count_28_io_out ? io_r_218_b : _GEN_11597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11599 = 9'hdb == r_count_28_io_out ? io_r_219_b : _GEN_11598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11600 = 9'hdc == r_count_28_io_out ? io_r_220_b : _GEN_11599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11601 = 9'hdd == r_count_28_io_out ? io_r_221_b : _GEN_11600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11602 = 9'hde == r_count_28_io_out ? io_r_222_b : _GEN_11601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11603 = 9'hdf == r_count_28_io_out ? io_r_223_b : _GEN_11602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11604 = 9'he0 == r_count_28_io_out ? io_r_224_b : _GEN_11603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11605 = 9'he1 == r_count_28_io_out ? io_r_225_b : _GEN_11604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11606 = 9'he2 == r_count_28_io_out ? io_r_226_b : _GEN_11605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11607 = 9'he3 == r_count_28_io_out ? io_r_227_b : _GEN_11606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11608 = 9'he4 == r_count_28_io_out ? io_r_228_b : _GEN_11607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11609 = 9'he5 == r_count_28_io_out ? io_r_229_b : _GEN_11608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11610 = 9'he6 == r_count_28_io_out ? io_r_230_b : _GEN_11609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11611 = 9'he7 == r_count_28_io_out ? io_r_231_b : _GEN_11610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11612 = 9'he8 == r_count_28_io_out ? io_r_232_b : _GEN_11611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11613 = 9'he9 == r_count_28_io_out ? io_r_233_b : _GEN_11612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11614 = 9'hea == r_count_28_io_out ? io_r_234_b : _GEN_11613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11615 = 9'heb == r_count_28_io_out ? io_r_235_b : _GEN_11614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11616 = 9'hec == r_count_28_io_out ? io_r_236_b : _GEN_11615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11617 = 9'hed == r_count_28_io_out ? io_r_237_b : _GEN_11616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11618 = 9'hee == r_count_28_io_out ? io_r_238_b : _GEN_11617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11619 = 9'hef == r_count_28_io_out ? io_r_239_b : _GEN_11618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11620 = 9'hf0 == r_count_28_io_out ? io_r_240_b : _GEN_11619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11621 = 9'hf1 == r_count_28_io_out ? io_r_241_b : _GEN_11620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11622 = 9'hf2 == r_count_28_io_out ? io_r_242_b : _GEN_11621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11623 = 9'hf3 == r_count_28_io_out ? io_r_243_b : _GEN_11622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11624 = 9'hf4 == r_count_28_io_out ? io_r_244_b : _GEN_11623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11625 = 9'hf5 == r_count_28_io_out ? io_r_245_b : _GEN_11624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11626 = 9'hf6 == r_count_28_io_out ? io_r_246_b : _GEN_11625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11627 = 9'hf7 == r_count_28_io_out ? io_r_247_b : _GEN_11626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11628 = 9'hf8 == r_count_28_io_out ? io_r_248_b : _GEN_11627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11629 = 9'hf9 == r_count_28_io_out ? io_r_249_b : _GEN_11628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11630 = 9'hfa == r_count_28_io_out ? io_r_250_b : _GEN_11629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11631 = 9'hfb == r_count_28_io_out ? io_r_251_b : _GEN_11630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11632 = 9'hfc == r_count_28_io_out ? io_r_252_b : _GEN_11631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11633 = 9'hfd == r_count_28_io_out ? io_r_253_b : _GEN_11632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11634 = 9'hfe == r_count_28_io_out ? io_r_254_b : _GEN_11633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11635 = 9'hff == r_count_28_io_out ? io_r_255_b : _GEN_11634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11636 = 9'h100 == r_count_28_io_out ? io_r_256_b : _GEN_11635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11637 = 9'h101 == r_count_28_io_out ? io_r_257_b : _GEN_11636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11638 = 9'h102 == r_count_28_io_out ? io_r_258_b : _GEN_11637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11639 = 9'h103 == r_count_28_io_out ? io_r_259_b : _GEN_11638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11640 = 9'h104 == r_count_28_io_out ? io_r_260_b : _GEN_11639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11641 = 9'h105 == r_count_28_io_out ? io_r_261_b : _GEN_11640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11642 = 9'h106 == r_count_28_io_out ? io_r_262_b : _GEN_11641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11643 = 9'h107 == r_count_28_io_out ? io_r_263_b : _GEN_11642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11644 = 9'h108 == r_count_28_io_out ? io_r_264_b : _GEN_11643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11645 = 9'h109 == r_count_28_io_out ? io_r_265_b : _GEN_11644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11646 = 9'h10a == r_count_28_io_out ? io_r_266_b : _GEN_11645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11647 = 9'h10b == r_count_28_io_out ? io_r_267_b : _GEN_11646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11648 = 9'h10c == r_count_28_io_out ? io_r_268_b : _GEN_11647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11649 = 9'h10d == r_count_28_io_out ? io_r_269_b : _GEN_11648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11650 = 9'h10e == r_count_28_io_out ? io_r_270_b : _GEN_11649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11651 = 9'h10f == r_count_28_io_out ? io_r_271_b : _GEN_11650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11652 = 9'h110 == r_count_28_io_out ? io_r_272_b : _GEN_11651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11653 = 9'h111 == r_count_28_io_out ? io_r_273_b : _GEN_11652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11654 = 9'h112 == r_count_28_io_out ? io_r_274_b : _GEN_11653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11655 = 9'h113 == r_count_28_io_out ? io_r_275_b : _GEN_11654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11656 = 9'h114 == r_count_28_io_out ? io_r_276_b : _GEN_11655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11657 = 9'h115 == r_count_28_io_out ? io_r_277_b : _GEN_11656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11658 = 9'h116 == r_count_28_io_out ? io_r_278_b : _GEN_11657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11659 = 9'h117 == r_count_28_io_out ? io_r_279_b : _GEN_11658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11660 = 9'h118 == r_count_28_io_out ? io_r_280_b : _GEN_11659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11661 = 9'h119 == r_count_28_io_out ? io_r_281_b : _GEN_11660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11662 = 9'h11a == r_count_28_io_out ? io_r_282_b : _GEN_11661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11663 = 9'h11b == r_count_28_io_out ? io_r_283_b : _GEN_11662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11664 = 9'h11c == r_count_28_io_out ? io_r_284_b : _GEN_11663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11665 = 9'h11d == r_count_28_io_out ? io_r_285_b : _GEN_11664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11666 = 9'h11e == r_count_28_io_out ? io_r_286_b : _GEN_11665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11667 = 9'h11f == r_count_28_io_out ? io_r_287_b : _GEN_11666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11668 = 9'h120 == r_count_28_io_out ? io_r_288_b : _GEN_11667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11669 = 9'h121 == r_count_28_io_out ? io_r_289_b : _GEN_11668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11670 = 9'h122 == r_count_28_io_out ? io_r_290_b : _GEN_11669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11671 = 9'h123 == r_count_28_io_out ? io_r_291_b : _GEN_11670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11672 = 9'h124 == r_count_28_io_out ? io_r_292_b : _GEN_11671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11673 = 9'h125 == r_count_28_io_out ? io_r_293_b : _GEN_11672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11674 = 9'h126 == r_count_28_io_out ? io_r_294_b : _GEN_11673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11675 = 9'h127 == r_count_28_io_out ? io_r_295_b : _GEN_11674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11676 = 9'h128 == r_count_28_io_out ? io_r_296_b : _GEN_11675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11677 = 9'h129 == r_count_28_io_out ? io_r_297_b : _GEN_11676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11678 = 9'h12a == r_count_28_io_out ? io_r_298_b : _GEN_11677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11679 = 9'h12b == r_count_28_io_out ? io_r_299_b : _GEN_11678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11680 = 9'h12c == r_count_28_io_out ? io_r_300_b : _GEN_11679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11681 = 9'h12d == r_count_28_io_out ? io_r_301_b : _GEN_11680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11682 = 9'h12e == r_count_28_io_out ? io_r_302_b : _GEN_11681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11683 = 9'h12f == r_count_28_io_out ? io_r_303_b : _GEN_11682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11684 = 9'h130 == r_count_28_io_out ? io_r_304_b : _GEN_11683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11685 = 9'h131 == r_count_28_io_out ? io_r_305_b : _GEN_11684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11686 = 9'h132 == r_count_28_io_out ? io_r_306_b : _GEN_11685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11687 = 9'h133 == r_count_28_io_out ? io_r_307_b : _GEN_11686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11688 = 9'h134 == r_count_28_io_out ? io_r_308_b : _GEN_11687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11689 = 9'h135 == r_count_28_io_out ? io_r_309_b : _GEN_11688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11690 = 9'h136 == r_count_28_io_out ? io_r_310_b : _GEN_11689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11691 = 9'h137 == r_count_28_io_out ? io_r_311_b : _GEN_11690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11692 = 9'h138 == r_count_28_io_out ? io_r_312_b : _GEN_11691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11693 = 9'h139 == r_count_28_io_out ? io_r_313_b : _GEN_11692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11694 = 9'h13a == r_count_28_io_out ? io_r_314_b : _GEN_11693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11695 = 9'h13b == r_count_28_io_out ? io_r_315_b : _GEN_11694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11696 = 9'h13c == r_count_28_io_out ? io_r_316_b : _GEN_11695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11697 = 9'h13d == r_count_28_io_out ? io_r_317_b : _GEN_11696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11698 = 9'h13e == r_count_28_io_out ? io_r_318_b : _GEN_11697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11699 = 9'h13f == r_count_28_io_out ? io_r_319_b : _GEN_11698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11700 = 9'h140 == r_count_28_io_out ? io_r_320_b : _GEN_11699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11701 = 9'h141 == r_count_28_io_out ? io_r_321_b : _GEN_11700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11702 = 9'h142 == r_count_28_io_out ? io_r_322_b : _GEN_11701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11703 = 9'h143 == r_count_28_io_out ? io_r_323_b : _GEN_11702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11704 = 9'h144 == r_count_28_io_out ? io_r_324_b : _GEN_11703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11705 = 9'h145 == r_count_28_io_out ? io_r_325_b : _GEN_11704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11706 = 9'h146 == r_count_28_io_out ? io_r_326_b : _GEN_11705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11707 = 9'h147 == r_count_28_io_out ? io_r_327_b : _GEN_11706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11708 = 9'h148 == r_count_28_io_out ? io_r_328_b : _GEN_11707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11709 = 9'h149 == r_count_28_io_out ? io_r_329_b : _GEN_11708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11710 = 9'h14a == r_count_28_io_out ? io_r_330_b : _GEN_11709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11711 = 9'h14b == r_count_28_io_out ? io_r_331_b : _GEN_11710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11712 = 9'h14c == r_count_28_io_out ? io_r_332_b : _GEN_11711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11713 = 9'h14d == r_count_28_io_out ? io_r_333_b : _GEN_11712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11714 = 9'h14e == r_count_28_io_out ? io_r_334_b : _GEN_11713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11715 = 9'h14f == r_count_28_io_out ? io_r_335_b : _GEN_11714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11716 = 9'h150 == r_count_28_io_out ? io_r_336_b : _GEN_11715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11717 = 9'h151 == r_count_28_io_out ? io_r_337_b : _GEN_11716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11718 = 9'h152 == r_count_28_io_out ? io_r_338_b : _GEN_11717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11719 = 9'h153 == r_count_28_io_out ? io_r_339_b : _GEN_11718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11720 = 9'h154 == r_count_28_io_out ? io_r_340_b : _GEN_11719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11721 = 9'h155 == r_count_28_io_out ? io_r_341_b : _GEN_11720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11722 = 9'h156 == r_count_28_io_out ? io_r_342_b : _GEN_11721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11723 = 9'h157 == r_count_28_io_out ? io_r_343_b : _GEN_11722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11724 = 9'h158 == r_count_28_io_out ? io_r_344_b : _GEN_11723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11725 = 9'h159 == r_count_28_io_out ? io_r_345_b : _GEN_11724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11726 = 9'h15a == r_count_28_io_out ? io_r_346_b : _GEN_11725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11727 = 9'h15b == r_count_28_io_out ? io_r_347_b : _GEN_11726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11728 = 9'h15c == r_count_28_io_out ? io_r_348_b : _GEN_11727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11729 = 9'h15d == r_count_28_io_out ? io_r_349_b : _GEN_11728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11730 = 9'h15e == r_count_28_io_out ? io_r_350_b : _GEN_11729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11731 = 9'h15f == r_count_28_io_out ? io_r_351_b : _GEN_11730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11732 = 9'h160 == r_count_28_io_out ? io_r_352_b : _GEN_11731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11733 = 9'h161 == r_count_28_io_out ? io_r_353_b : _GEN_11732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11734 = 9'h162 == r_count_28_io_out ? io_r_354_b : _GEN_11733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11735 = 9'h163 == r_count_28_io_out ? io_r_355_b : _GEN_11734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11736 = 9'h164 == r_count_28_io_out ? io_r_356_b : _GEN_11735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11737 = 9'h165 == r_count_28_io_out ? io_r_357_b : _GEN_11736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11738 = 9'h166 == r_count_28_io_out ? io_r_358_b : _GEN_11737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11739 = 9'h167 == r_count_28_io_out ? io_r_359_b : _GEN_11738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11740 = 9'h168 == r_count_28_io_out ? io_r_360_b : _GEN_11739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11741 = 9'h169 == r_count_28_io_out ? io_r_361_b : _GEN_11740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11742 = 9'h16a == r_count_28_io_out ? io_r_362_b : _GEN_11741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11743 = 9'h16b == r_count_28_io_out ? io_r_363_b : _GEN_11742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11744 = 9'h16c == r_count_28_io_out ? io_r_364_b : _GEN_11743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11745 = 9'h16d == r_count_28_io_out ? io_r_365_b : _GEN_11744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11746 = 9'h16e == r_count_28_io_out ? io_r_366_b : _GEN_11745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11747 = 9'h16f == r_count_28_io_out ? io_r_367_b : _GEN_11746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11748 = 9'h170 == r_count_28_io_out ? io_r_368_b : _GEN_11747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11749 = 9'h171 == r_count_28_io_out ? io_r_369_b : _GEN_11748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11750 = 9'h172 == r_count_28_io_out ? io_r_370_b : _GEN_11749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11751 = 9'h173 == r_count_28_io_out ? io_r_371_b : _GEN_11750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11752 = 9'h174 == r_count_28_io_out ? io_r_372_b : _GEN_11751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11753 = 9'h175 == r_count_28_io_out ? io_r_373_b : _GEN_11752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11754 = 9'h176 == r_count_28_io_out ? io_r_374_b : _GEN_11753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11755 = 9'h177 == r_count_28_io_out ? io_r_375_b : _GEN_11754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11756 = 9'h178 == r_count_28_io_out ? io_r_376_b : _GEN_11755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11757 = 9'h179 == r_count_28_io_out ? io_r_377_b : _GEN_11756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11758 = 9'h17a == r_count_28_io_out ? io_r_378_b : _GEN_11757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11759 = 9'h17b == r_count_28_io_out ? io_r_379_b : _GEN_11758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11760 = 9'h17c == r_count_28_io_out ? io_r_380_b : _GEN_11759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11761 = 9'h17d == r_count_28_io_out ? io_r_381_b : _GEN_11760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11762 = 9'h17e == r_count_28_io_out ? io_r_382_b : _GEN_11761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11763 = 9'h17f == r_count_28_io_out ? io_r_383_b : _GEN_11762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11764 = 9'h180 == r_count_28_io_out ? io_r_384_b : _GEN_11763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11765 = 9'h181 == r_count_28_io_out ? io_r_385_b : _GEN_11764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11766 = 9'h182 == r_count_28_io_out ? io_r_386_b : _GEN_11765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11767 = 9'h183 == r_count_28_io_out ? io_r_387_b : _GEN_11766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11768 = 9'h184 == r_count_28_io_out ? io_r_388_b : _GEN_11767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11769 = 9'h185 == r_count_28_io_out ? io_r_389_b : _GEN_11768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11770 = 9'h186 == r_count_28_io_out ? io_r_390_b : _GEN_11769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11771 = 9'h187 == r_count_28_io_out ? io_r_391_b : _GEN_11770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11772 = 9'h188 == r_count_28_io_out ? io_r_392_b : _GEN_11771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11773 = 9'h189 == r_count_28_io_out ? io_r_393_b : _GEN_11772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11774 = 9'h18a == r_count_28_io_out ? io_r_394_b : _GEN_11773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11775 = 9'h18b == r_count_28_io_out ? io_r_395_b : _GEN_11774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11776 = 9'h18c == r_count_28_io_out ? io_r_396_b : _GEN_11775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11777 = 9'h18d == r_count_28_io_out ? io_r_397_b : _GEN_11776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11778 = 9'h18e == r_count_28_io_out ? io_r_398_b : _GEN_11777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11781 = 9'h1 == r_count_29_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11782 = 9'h2 == r_count_29_io_out ? io_r_2_b : _GEN_11781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11783 = 9'h3 == r_count_29_io_out ? io_r_3_b : _GEN_11782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11784 = 9'h4 == r_count_29_io_out ? io_r_4_b : _GEN_11783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11785 = 9'h5 == r_count_29_io_out ? io_r_5_b : _GEN_11784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11786 = 9'h6 == r_count_29_io_out ? io_r_6_b : _GEN_11785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11787 = 9'h7 == r_count_29_io_out ? io_r_7_b : _GEN_11786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11788 = 9'h8 == r_count_29_io_out ? io_r_8_b : _GEN_11787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11789 = 9'h9 == r_count_29_io_out ? io_r_9_b : _GEN_11788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11790 = 9'ha == r_count_29_io_out ? io_r_10_b : _GEN_11789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11791 = 9'hb == r_count_29_io_out ? io_r_11_b : _GEN_11790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11792 = 9'hc == r_count_29_io_out ? io_r_12_b : _GEN_11791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11793 = 9'hd == r_count_29_io_out ? io_r_13_b : _GEN_11792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11794 = 9'he == r_count_29_io_out ? io_r_14_b : _GEN_11793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11795 = 9'hf == r_count_29_io_out ? io_r_15_b : _GEN_11794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11796 = 9'h10 == r_count_29_io_out ? io_r_16_b : _GEN_11795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11797 = 9'h11 == r_count_29_io_out ? io_r_17_b : _GEN_11796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11798 = 9'h12 == r_count_29_io_out ? io_r_18_b : _GEN_11797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11799 = 9'h13 == r_count_29_io_out ? io_r_19_b : _GEN_11798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11800 = 9'h14 == r_count_29_io_out ? io_r_20_b : _GEN_11799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11801 = 9'h15 == r_count_29_io_out ? io_r_21_b : _GEN_11800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11802 = 9'h16 == r_count_29_io_out ? io_r_22_b : _GEN_11801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11803 = 9'h17 == r_count_29_io_out ? io_r_23_b : _GEN_11802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11804 = 9'h18 == r_count_29_io_out ? io_r_24_b : _GEN_11803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11805 = 9'h19 == r_count_29_io_out ? io_r_25_b : _GEN_11804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11806 = 9'h1a == r_count_29_io_out ? io_r_26_b : _GEN_11805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11807 = 9'h1b == r_count_29_io_out ? io_r_27_b : _GEN_11806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11808 = 9'h1c == r_count_29_io_out ? io_r_28_b : _GEN_11807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11809 = 9'h1d == r_count_29_io_out ? io_r_29_b : _GEN_11808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11810 = 9'h1e == r_count_29_io_out ? io_r_30_b : _GEN_11809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11811 = 9'h1f == r_count_29_io_out ? io_r_31_b : _GEN_11810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11812 = 9'h20 == r_count_29_io_out ? io_r_32_b : _GEN_11811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11813 = 9'h21 == r_count_29_io_out ? io_r_33_b : _GEN_11812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11814 = 9'h22 == r_count_29_io_out ? io_r_34_b : _GEN_11813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11815 = 9'h23 == r_count_29_io_out ? io_r_35_b : _GEN_11814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11816 = 9'h24 == r_count_29_io_out ? io_r_36_b : _GEN_11815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11817 = 9'h25 == r_count_29_io_out ? io_r_37_b : _GEN_11816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11818 = 9'h26 == r_count_29_io_out ? io_r_38_b : _GEN_11817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11819 = 9'h27 == r_count_29_io_out ? io_r_39_b : _GEN_11818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11820 = 9'h28 == r_count_29_io_out ? io_r_40_b : _GEN_11819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11821 = 9'h29 == r_count_29_io_out ? io_r_41_b : _GEN_11820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11822 = 9'h2a == r_count_29_io_out ? io_r_42_b : _GEN_11821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11823 = 9'h2b == r_count_29_io_out ? io_r_43_b : _GEN_11822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11824 = 9'h2c == r_count_29_io_out ? io_r_44_b : _GEN_11823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11825 = 9'h2d == r_count_29_io_out ? io_r_45_b : _GEN_11824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11826 = 9'h2e == r_count_29_io_out ? io_r_46_b : _GEN_11825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11827 = 9'h2f == r_count_29_io_out ? io_r_47_b : _GEN_11826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11828 = 9'h30 == r_count_29_io_out ? io_r_48_b : _GEN_11827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11829 = 9'h31 == r_count_29_io_out ? io_r_49_b : _GEN_11828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11830 = 9'h32 == r_count_29_io_out ? io_r_50_b : _GEN_11829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11831 = 9'h33 == r_count_29_io_out ? io_r_51_b : _GEN_11830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11832 = 9'h34 == r_count_29_io_out ? io_r_52_b : _GEN_11831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11833 = 9'h35 == r_count_29_io_out ? io_r_53_b : _GEN_11832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11834 = 9'h36 == r_count_29_io_out ? io_r_54_b : _GEN_11833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11835 = 9'h37 == r_count_29_io_out ? io_r_55_b : _GEN_11834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11836 = 9'h38 == r_count_29_io_out ? io_r_56_b : _GEN_11835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11837 = 9'h39 == r_count_29_io_out ? io_r_57_b : _GEN_11836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11838 = 9'h3a == r_count_29_io_out ? io_r_58_b : _GEN_11837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11839 = 9'h3b == r_count_29_io_out ? io_r_59_b : _GEN_11838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11840 = 9'h3c == r_count_29_io_out ? io_r_60_b : _GEN_11839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11841 = 9'h3d == r_count_29_io_out ? io_r_61_b : _GEN_11840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11842 = 9'h3e == r_count_29_io_out ? io_r_62_b : _GEN_11841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11843 = 9'h3f == r_count_29_io_out ? io_r_63_b : _GEN_11842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11844 = 9'h40 == r_count_29_io_out ? io_r_64_b : _GEN_11843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11845 = 9'h41 == r_count_29_io_out ? io_r_65_b : _GEN_11844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11846 = 9'h42 == r_count_29_io_out ? io_r_66_b : _GEN_11845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11847 = 9'h43 == r_count_29_io_out ? io_r_67_b : _GEN_11846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11848 = 9'h44 == r_count_29_io_out ? io_r_68_b : _GEN_11847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11849 = 9'h45 == r_count_29_io_out ? io_r_69_b : _GEN_11848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11850 = 9'h46 == r_count_29_io_out ? io_r_70_b : _GEN_11849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11851 = 9'h47 == r_count_29_io_out ? io_r_71_b : _GEN_11850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11852 = 9'h48 == r_count_29_io_out ? io_r_72_b : _GEN_11851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11853 = 9'h49 == r_count_29_io_out ? io_r_73_b : _GEN_11852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11854 = 9'h4a == r_count_29_io_out ? io_r_74_b : _GEN_11853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11855 = 9'h4b == r_count_29_io_out ? io_r_75_b : _GEN_11854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11856 = 9'h4c == r_count_29_io_out ? io_r_76_b : _GEN_11855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11857 = 9'h4d == r_count_29_io_out ? io_r_77_b : _GEN_11856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11858 = 9'h4e == r_count_29_io_out ? io_r_78_b : _GEN_11857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11859 = 9'h4f == r_count_29_io_out ? io_r_79_b : _GEN_11858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11860 = 9'h50 == r_count_29_io_out ? io_r_80_b : _GEN_11859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11861 = 9'h51 == r_count_29_io_out ? io_r_81_b : _GEN_11860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11862 = 9'h52 == r_count_29_io_out ? io_r_82_b : _GEN_11861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11863 = 9'h53 == r_count_29_io_out ? io_r_83_b : _GEN_11862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11864 = 9'h54 == r_count_29_io_out ? io_r_84_b : _GEN_11863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11865 = 9'h55 == r_count_29_io_out ? io_r_85_b : _GEN_11864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11866 = 9'h56 == r_count_29_io_out ? io_r_86_b : _GEN_11865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11867 = 9'h57 == r_count_29_io_out ? io_r_87_b : _GEN_11866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11868 = 9'h58 == r_count_29_io_out ? io_r_88_b : _GEN_11867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11869 = 9'h59 == r_count_29_io_out ? io_r_89_b : _GEN_11868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11870 = 9'h5a == r_count_29_io_out ? io_r_90_b : _GEN_11869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11871 = 9'h5b == r_count_29_io_out ? io_r_91_b : _GEN_11870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11872 = 9'h5c == r_count_29_io_out ? io_r_92_b : _GEN_11871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11873 = 9'h5d == r_count_29_io_out ? io_r_93_b : _GEN_11872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11874 = 9'h5e == r_count_29_io_out ? io_r_94_b : _GEN_11873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11875 = 9'h5f == r_count_29_io_out ? io_r_95_b : _GEN_11874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11876 = 9'h60 == r_count_29_io_out ? io_r_96_b : _GEN_11875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11877 = 9'h61 == r_count_29_io_out ? io_r_97_b : _GEN_11876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11878 = 9'h62 == r_count_29_io_out ? io_r_98_b : _GEN_11877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11879 = 9'h63 == r_count_29_io_out ? io_r_99_b : _GEN_11878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11880 = 9'h64 == r_count_29_io_out ? io_r_100_b : _GEN_11879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11881 = 9'h65 == r_count_29_io_out ? io_r_101_b : _GEN_11880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11882 = 9'h66 == r_count_29_io_out ? io_r_102_b : _GEN_11881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11883 = 9'h67 == r_count_29_io_out ? io_r_103_b : _GEN_11882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11884 = 9'h68 == r_count_29_io_out ? io_r_104_b : _GEN_11883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11885 = 9'h69 == r_count_29_io_out ? io_r_105_b : _GEN_11884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11886 = 9'h6a == r_count_29_io_out ? io_r_106_b : _GEN_11885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11887 = 9'h6b == r_count_29_io_out ? io_r_107_b : _GEN_11886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11888 = 9'h6c == r_count_29_io_out ? io_r_108_b : _GEN_11887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11889 = 9'h6d == r_count_29_io_out ? io_r_109_b : _GEN_11888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11890 = 9'h6e == r_count_29_io_out ? io_r_110_b : _GEN_11889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11891 = 9'h6f == r_count_29_io_out ? io_r_111_b : _GEN_11890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11892 = 9'h70 == r_count_29_io_out ? io_r_112_b : _GEN_11891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11893 = 9'h71 == r_count_29_io_out ? io_r_113_b : _GEN_11892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11894 = 9'h72 == r_count_29_io_out ? io_r_114_b : _GEN_11893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11895 = 9'h73 == r_count_29_io_out ? io_r_115_b : _GEN_11894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11896 = 9'h74 == r_count_29_io_out ? io_r_116_b : _GEN_11895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11897 = 9'h75 == r_count_29_io_out ? io_r_117_b : _GEN_11896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11898 = 9'h76 == r_count_29_io_out ? io_r_118_b : _GEN_11897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11899 = 9'h77 == r_count_29_io_out ? io_r_119_b : _GEN_11898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11900 = 9'h78 == r_count_29_io_out ? io_r_120_b : _GEN_11899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11901 = 9'h79 == r_count_29_io_out ? io_r_121_b : _GEN_11900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11902 = 9'h7a == r_count_29_io_out ? io_r_122_b : _GEN_11901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11903 = 9'h7b == r_count_29_io_out ? io_r_123_b : _GEN_11902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11904 = 9'h7c == r_count_29_io_out ? io_r_124_b : _GEN_11903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11905 = 9'h7d == r_count_29_io_out ? io_r_125_b : _GEN_11904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11906 = 9'h7e == r_count_29_io_out ? io_r_126_b : _GEN_11905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11907 = 9'h7f == r_count_29_io_out ? io_r_127_b : _GEN_11906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11908 = 9'h80 == r_count_29_io_out ? io_r_128_b : _GEN_11907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11909 = 9'h81 == r_count_29_io_out ? io_r_129_b : _GEN_11908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11910 = 9'h82 == r_count_29_io_out ? io_r_130_b : _GEN_11909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11911 = 9'h83 == r_count_29_io_out ? io_r_131_b : _GEN_11910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11912 = 9'h84 == r_count_29_io_out ? io_r_132_b : _GEN_11911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11913 = 9'h85 == r_count_29_io_out ? io_r_133_b : _GEN_11912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11914 = 9'h86 == r_count_29_io_out ? io_r_134_b : _GEN_11913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11915 = 9'h87 == r_count_29_io_out ? io_r_135_b : _GEN_11914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11916 = 9'h88 == r_count_29_io_out ? io_r_136_b : _GEN_11915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11917 = 9'h89 == r_count_29_io_out ? io_r_137_b : _GEN_11916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11918 = 9'h8a == r_count_29_io_out ? io_r_138_b : _GEN_11917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11919 = 9'h8b == r_count_29_io_out ? io_r_139_b : _GEN_11918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11920 = 9'h8c == r_count_29_io_out ? io_r_140_b : _GEN_11919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11921 = 9'h8d == r_count_29_io_out ? io_r_141_b : _GEN_11920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11922 = 9'h8e == r_count_29_io_out ? io_r_142_b : _GEN_11921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11923 = 9'h8f == r_count_29_io_out ? io_r_143_b : _GEN_11922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11924 = 9'h90 == r_count_29_io_out ? io_r_144_b : _GEN_11923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11925 = 9'h91 == r_count_29_io_out ? io_r_145_b : _GEN_11924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11926 = 9'h92 == r_count_29_io_out ? io_r_146_b : _GEN_11925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11927 = 9'h93 == r_count_29_io_out ? io_r_147_b : _GEN_11926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11928 = 9'h94 == r_count_29_io_out ? io_r_148_b : _GEN_11927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11929 = 9'h95 == r_count_29_io_out ? io_r_149_b : _GEN_11928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11930 = 9'h96 == r_count_29_io_out ? io_r_150_b : _GEN_11929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11931 = 9'h97 == r_count_29_io_out ? io_r_151_b : _GEN_11930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11932 = 9'h98 == r_count_29_io_out ? io_r_152_b : _GEN_11931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11933 = 9'h99 == r_count_29_io_out ? io_r_153_b : _GEN_11932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11934 = 9'h9a == r_count_29_io_out ? io_r_154_b : _GEN_11933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11935 = 9'h9b == r_count_29_io_out ? io_r_155_b : _GEN_11934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11936 = 9'h9c == r_count_29_io_out ? io_r_156_b : _GEN_11935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11937 = 9'h9d == r_count_29_io_out ? io_r_157_b : _GEN_11936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11938 = 9'h9e == r_count_29_io_out ? io_r_158_b : _GEN_11937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11939 = 9'h9f == r_count_29_io_out ? io_r_159_b : _GEN_11938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11940 = 9'ha0 == r_count_29_io_out ? io_r_160_b : _GEN_11939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11941 = 9'ha1 == r_count_29_io_out ? io_r_161_b : _GEN_11940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11942 = 9'ha2 == r_count_29_io_out ? io_r_162_b : _GEN_11941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11943 = 9'ha3 == r_count_29_io_out ? io_r_163_b : _GEN_11942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11944 = 9'ha4 == r_count_29_io_out ? io_r_164_b : _GEN_11943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11945 = 9'ha5 == r_count_29_io_out ? io_r_165_b : _GEN_11944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11946 = 9'ha6 == r_count_29_io_out ? io_r_166_b : _GEN_11945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11947 = 9'ha7 == r_count_29_io_out ? io_r_167_b : _GEN_11946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11948 = 9'ha8 == r_count_29_io_out ? io_r_168_b : _GEN_11947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11949 = 9'ha9 == r_count_29_io_out ? io_r_169_b : _GEN_11948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11950 = 9'haa == r_count_29_io_out ? io_r_170_b : _GEN_11949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11951 = 9'hab == r_count_29_io_out ? io_r_171_b : _GEN_11950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11952 = 9'hac == r_count_29_io_out ? io_r_172_b : _GEN_11951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11953 = 9'had == r_count_29_io_out ? io_r_173_b : _GEN_11952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11954 = 9'hae == r_count_29_io_out ? io_r_174_b : _GEN_11953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11955 = 9'haf == r_count_29_io_out ? io_r_175_b : _GEN_11954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11956 = 9'hb0 == r_count_29_io_out ? io_r_176_b : _GEN_11955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11957 = 9'hb1 == r_count_29_io_out ? io_r_177_b : _GEN_11956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11958 = 9'hb2 == r_count_29_io_out ? io_r_178_b : _GEN_11957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11959 = 9'hb3 == r_count_29_io_out ? io_r_179_b : _GEN_11958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11960 = 9'hb4 == r_count_29_io_out ? io_r_180_b : _GEN_11959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11961 = 9'hb5 == r_count_29_io_out ? io_r_181_b : _GEN_11960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11962 = 9'hb6 == r_count_29_io_out ? io_r_182_b : _GEN_11961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11963 = 9'hb7 == r_count_29_io_out ? io_r_183_b : _GEN_11962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11964 = 9'hb8 == r_count_29_io_out ? io_r_184_b : _GEN_11963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11965 = 9'hb9 == r_count_29_io_out ? io_r_185_b : _GEN_11964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11966 = 9'hba == r_count_29_io_out ? io_r_186_b : _GEN_11965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11967 = 9'hbb == r_count_29_io_out ? io_r_187_b : _GEN_11966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11968 = 9'hbc == r_count_29_io_out ? io_r_188_b : _GEN_11967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11969 = 9'hbd == r_count_29_io_out ? io_r_189_b : _GEN_11968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11970 = 9'hbe == r_count_29_io_out ? io_r_190_b : _GEN_11969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11971 = 9'hbf == r_count_29_io_out ? io_r_191_b : _GEN_11970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11972 = 9'hc0 == r_count_29_io_out ? io_r_192_b : _GEN_11971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11973 = 9'hc1 == r_count_29_io_out ? io_r_193_b : _GEN_11972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11974 = 9'hc2 == r_count_29_io_out ? io_r_194_b : _GEN_11973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11975 = 9'hc3 == r_count_29_io_out ? io_r_195_b : _GEN_11974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11976 = 9'hc4 == r_count_29_io_out ? io_r_196_b : _GEN_11975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11977 = 9'hc5 == r_count_29_io_out ? io_r_197_b : _GEN_11976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11978 = 9'hc6 == r_count_29_io_out ? io_r_198_b : _GEN_11977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11979 = 9'hc7 == r_count_29_io_out ? io_r_199_b : _GEN_11978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11980 = 9'hc8 == r_count_29_io_out ? io_r_200_b : _GEN_11979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11981 = 9'hc9 == r_count_29_io_out ? io_r_201_b : _GEN_11980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11982 = 9'hca == r_count_29_io_out ? io_r_202_b : _GEN_11981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11983 = 9'hcb == r_count_29_io_out ? io_r_203_b : _GEN_11982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11984 = 9'hcc == r_count_29_io_out ? io_r_204_b : _GEN_11983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11985 = 9'hcd == r_count_29_io_out ? io_r_205_b : _GEN_11984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11986 = 9'hce == r_count_29_io_out ? io_r_206_b : _GEN_11985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11987 = 9'hcf == r_count_29_io_out ? io_r_207_b : _GEN_11986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11988 = 9'hd0 == r_count_29_io_out ? io_r_208_b : _GEN_11987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11989 = 9'hd1 == r_count_29_io_out ? io_r_209_b : _GEN_11988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11990 = 9'hd2 == r_count_29_io_out ? io_r_210_b : _GEN_11989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11991 = 9'hd3 == r_count_29_io_out ? io_r_211_b : _GEN_11990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11992 = 9'hd4 == r_count_29_io_out ? io_r_212_b : _GEN_11991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11993 = 9'hd5 == r_count_29_io_out ? io_r_213_b : _GEN_11992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11994 = 9'hd6 == r_count_29_io_out ? io_r_214_b : _GEN_11993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11995 = 9'hd7 == r_count_29_io_out ? io_r_215_b : _GEN_11994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11996 = 9'hd8 == r_count_29_io_out ? io_r_216_b : _GEN_11995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11997 = 9'hd9 == r_count_29_io_out ? io_r_217_b : _GEN_11996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11998 = 9'hda == r_count_29_io_out ? io_r_218_b : _GEN_11997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11999 = 9'hdb == r_count_29_io_out ? io_r_219_b : _GEN_11998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12000 = 9'hdc == r_count_29_io_out ? io_r_220_b : _GEN_11999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12001 = 9'hdd == r_count_29_io_out ? io_r_221_b : _GEN_12000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12002 = 9'hde == r_count_29_io_out ? io_r_222_b : _GEN_12001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12003 = 9'hdf == r_count_29_io_out ? io_r_223_b : _GEN_12002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12004 = 9'he0 == r_count_29_io_out ? io_r_224_b : _GEN_12003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12005 = 9'he1 == r_count_29_io_out ? io_r_225_b : _GEN_12004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12006 = 9'he2 == r_count_29_io_out ? io_r_226_b : _GEN_12005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12007 = 9'he3 == r_count_29_io_out ? io_r_227_b : _GEN_12006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12008 = 9'he4 == r_count_29_io_out ? io_r_228_b : _GEN_12007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12009 = 9'he5 == r_count_29_io_out ? io_r_229_b : _GEN_12008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12010 = 9'he6 == r_count_29_io_out ? io_r_230_b : _GEN_12009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12011 = 9'he7 == r_count_29_io_out ? io_r_231_b : _GEN_12010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12012 = 9'he8 == r_count_29_io_out ? io_r_232_b : _GEN_12011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12013 = 9'he9 == r_count_29_io_out ? io_r_233_b : _GEN_12012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12014 = 9'hea == r_count_29_io_out ? io_r_234_b : _GEN_12013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12015 = 9'heb == r_count_29_io_out ? io_r_235_b : _GEN_12014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12016 = 9'hec == r_count_29_io_out ? io_r_236_b : _GEN_12015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12017 = 9'hed == r_count_29_io_out ? io_r_237_b : _GEN_12016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12018 = 9'hee == r_count_29_io_out ? io_r_238_b : _GEN_12017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12019 = 9'hef == r_count_29_io_out ? io_r_239_b : _GEN_12018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12020 = 9'hf0 == r_count_29_io_out ? io_r_240_b : _GEN_12019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12021 = 9'hf1 == r_count_29_io_out ? io_r_241_b : _GEN_12020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12022 = 9'hf2 == r_count_29_io_out ? io_r_242_b : _GEN_12021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12023 = 9'hf3 == r_count_29_io_out ? io_r_243_b : _GEN_12022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12024 = 9'hf4 == r_count_29_io_out ? io_r_244_b : _GEN_12023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12025 = 9'hf5 == r_count_29_io_out ? io_r_245_b : _GEN_12024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12026 = 9'hf6 == r_count_29_io_out ? io_r_246_b : _GEN_12025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12027 = 9'hf7 == r_count_29_io_out ? io_r_247_b : _GEN_12026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12028 = 9'hf8 == r_count_29_io_out ? io_r_248_b : _GEN_12027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12029 = 9'hf9 == r_count_29_io_out ? io_r_249_b : _GEN_12028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12030 = 9'hfa == r_count_29_io_out ? io_r_250_b : _GEN_12029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12031 = 9'hfb == r_count_29_io_out ? io_r_251_b : _GEN_12030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12032 = 9'hfc == r_count_29_io_out ? io_r_252_b : _GEN_12031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12033 = 9'hfd == r_count_29_io_out ? io_r_253_b : _GEN_12032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12034 = 9'hfe == r_count_29_io_out ? io_r_254_b : _GEN_12033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12035 = 9'hff == r_count_29_io_out ? io_r_255_b : _GEN_12034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12036 = 9'h100 == r_count_29_io_out ? io_r_256_b : _GEN_12035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12037 = 9'h101 == r_count_29_io_out ? io_r_257_b : _GEN_12036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12038 = 9'h102 == r_count_29_io_out ? io_r_258_b : _GEN_12037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12039 = 9'h103 == r_count_29_io_out ? io_r_259_b : _GEN_12038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12040 = 9'h104 == r_count_29_io_out ? io_r_260_b : _GEN_12039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12041 = 9'h105 == r_count_29_io_out ? io_r_261_b : _GEN_12040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12042 = 9'h106 == r_count_29_io_out ? io_r_262_b : _GEN_12041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12043 = 9'h107 == r_count_29_io_out ? io_r_263_b : _GEN_12042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12044 = 9'h108 == r_count_29_io_out ? io_r_264_b : _GEN_12043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12045 = 9'h109 == r_count_29_io_out ? io_r_265_b : _GEN_12044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12046 = 9'h10a == r_count_29_io_out ? io_r_266_b : _GEN_12045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12047 = 9'h10b == r_count_29_io_out ? io_r_267_b : _GEN_12046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12048 = 9'h10c == r_count_29_io_out ? io_r_268_b : _GEN_12047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12049 = 9'h10d == r_count_29_io_out ? io_r_269_b : _GEN_12048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12050 = 9'h10e == r_count_29_io_out ? io_r_270_b : _GEN_12049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12051 = 9'h10f == r_count_29_io_out ? io_r_271_b : _GEN_12050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12052 = 9'h110 == r_count_29_io_out ? io_r_272_b : _GEN_12051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12053 = 9'h111 == r_count_29_io_out ? io_r_273_b : _GEN_12052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12054 = 9'h112 == r_count_29_io_out ? io_r_274_b : _GEN_12053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12055 = 9'h113 == r_count_29_io_out ? io_r_275_b : _GEN_12054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12056 = 9'h114 == r_count_29_io_out ? io_r_276_b : _GEN_12055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12057 = 9'h115 == r_count_29_io_out ? io_r_277_b : _GEN_12056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12058 = 9'h116 == r_count_29_io_out ? io_r_278_b : _GEN_12057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12059 = 9'h117 == r_count_29_io_out ? io_r_279_b : _GEN_12058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12060 = 9'h118 == r_count_29_io_out ? io_r_280_b : _GEN_12059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12061 = 9'h119 == r_count_29_io_out ? io_r_281_b : _GEN_12060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12062 = 9'h11a == r_count_29_io_out ? io_r_282_b : _GEN_12061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12063 = 9'h11b == r_count_29_io_out ? io_r_283_b : _GEN_12062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12064 = 9'h11c == r_count_29_io_out ? io_r_284_b : _GEN_12063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12065 = 9'h11d == r_count_29_io_out ? io_r_285_b : _GEN_12064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12066 = 9'h11e == r_count_29_io_out ? io_r_286_b : _GEN_12065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12067 = 9'h11f == r_count_29_io_out ? io_r_287_b : _GEN_12066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12068 = 9'h120 == r_count_29_io_out ? io_r_288_b : _GEN_12067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12069 = 9'h121 == r_count_29_io_out ? io_r_289_b : _GEN_12068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12070 = 9'h122 == r_count_29_io_out ? io_r_290_b : _GEN_12069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12071 = 9'h123 == r_count_29_io_out ? io_r_291_b : _GEN_12070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12072 = 9'h124 == r_count_29_io_out ? io_r_292_b : _GEN_12071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12073 = 9'h125 == r_count_29_io_out ? io_r_293_b : _GEN_12072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12074 = 9'h126 == r_count_29_io_out ? io_r_294_b : _GEN_12073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12075 = 9'h127 == r_count_29_io_out ? io_r_295_b : _GEN_12074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12076 = 9'h128 == r_count_29_io_out ? io_r_296_b : _GEN_12075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12077 = 9'h129 == r_count_29_io_out ? io_r_297_b : _GEN_12076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12078 = 9'h12a == r_count_29_io_out ? io_r_298_b : _GEN_12077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12079 = 9'h12b == r_count_29_io_out ? io_r_299_b : _GEN_12078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12080 = 9'h12c == r_count_29_io_out ? io_r_300_b : _GEN_12079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12081 = 9'h12d == r_count_29_io_out ? io_r_301_b : _GEN_12080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12082 = 9'h12e == r_count_29_io_out ? io_r_302_b : _GEN_12081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12083 = 9'h12f == r_count_29_io_out ? io_r_303_b : _GEN_12082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12084 = 9'h130 == r_count_29_io_out ? io_r_304_b : _GEN_12083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12085 = 9'h131 == r_count_29_io_out ? io_r_305_b : _GEN_12084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12086 = 9'h132 == r_count_29_io_out ? io_r_306_b : _GEN_12085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12087 = 9'h133 == r_count_29_io_out ? io_r_307_b : _GEN_12086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12088 = 9'h134 == r_count_29_io_out ? io_r_308_b : _GEN_12087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12089 = 9'h135 == r_count_29_io_out ? io_r_309_b : _GEN_12088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12090 = 9'h136 == r_count_29_io_out ? io_r_310_b : _GEN_12089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12091 = 9'h137 == r_count_29_io_out ? io_r_311_b : _GEN_12090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12092 = 9'h138 == r_count_29_io_out ? io_r_312_b : _GEN_12091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12093 = 9'h139 == r_count_29_io_out ? io_r_313_b : _GEN_12092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12094 = 9'h13a == r_count_29_io_out ? io_r_314_b : _GEN_12093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12095 = 9'h13b == r_count_29_io_out ? io_r_315_b : _GEN_12094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12096 = 9'h13c == r_count_29_io_out ? io_r_316_b : _GEN_12095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12097 = 9'h13d == r_count_29_io_out ? io_r_317_b : _GEN_12096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12098 = 9'h13e == r_count_29_io_out ? io_r_318_b : _GEN_12097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12099 = 9'h13f == r_count_29_io_out ? io_r_319_b : _GEN_12098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12100 = 9'h140 == r_count_29_io_out ? io_r_320_b : _GEN_12099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12101 = 9'h141 == r_count_29_io_out ? io_r_321_b : _GEN_12100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12102 = 9'h142 == r_count_29_io_out ? io_r_322_b : _GEN_12101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12103 = 9'h143 == r_count_29_io_out ? io_r_323_b : _GEN_12102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12104 = 9'h144 == r_count_29_io_out ? io_r_324_b : _GEN_12103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12105 = 9'h145 == r_count_29_io_out ? io_r_325_b : _GEN_12104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12106 = 9'h146 == r_count_29_io_out ? io_r_326_b : _GEN_12105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12107 = 9'h147 == r_count_29_io_out ? io_r_327_b : _GEN_12106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12108 = 9'h148 == r_count_29_io_out ? io_r_328_b : _GEN_12107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12109 = 9'h149 == r_count_29_io_out ? io_r_329_b : _GEN_12108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12110 = 9'h14a == r_count_29_io_out ? io_r_330_b : _GEN_12109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12111 = 9'h14b == r_count_29_io_out ? io_r_331_b : _GEN_12110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12112 = 9'h14c == r_count_29_io_out ? io_r_332_b : _GEN_12111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12113 = 9'h14d == r_count_29_io_out ? io_r_333_b : _GEN_12112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12114 = 9'h14e == r_count_29_io_out ? io_r_334_b : _GEN_12113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12115 = 9'h14f == r_count_29_io_out ? io_r_335_b : _GEN_12114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12116 = 9'h150 == r_count_29_io_out ? io_r_336_b : _GEN_12115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12117 = 9'h151 == r_count_29_io_out ? io_r_337_b : _GEN_12116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12118 = 9'h152 == r_count_29_io_out ? io_r_338_b : _GEN_12117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12119 = 9'h153 == r_count_29_io_out ? io_r_339_b : _GEN_12118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12120 = 9'h154 == r_count_29_io_out ? io_r_340_b : _GEN_12119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12121 = 9'h155 == r_count_29_io_out ? io_r_341_b : _GEN_12120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12122 = 9'h156 == r_count_29_io_out ? io_r_342_b : _GEN_12121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12123 = 9'h157 == r_count_29_io_out ? io_r_343_b : _GEN_12122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12124 = 9'h158 == r_count_29_io_out ? io_r_344_b : _GEN_12123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12125 = 9'h159 == r_count_29_io_out ? io_r_345_b : _GEN_12124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12126 = 9'h15a == r_count_29_io_out ? io_r_346_b : _GEN_12125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12127 = 9'h15b == r_count_29_io_out ? io_r_347_b : _GEN_12126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12128 = 9'h15c == r_count_29_io_out ? io_r_348_b : _GEN_12127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12129 = 9'h15d == r_count_29_io_out ? io_r_349_b : _GEN_12128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12130 = 9'h15e == r_count_29_io_out ? io_r_350_b : _GEN_12129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12131 = 9'h15f == r_count_29_io_out ? io_r_351_b : _GEN_12130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12132 = 9'h160 == r_count_29_io_out ? io_r_352_b : _GEN_12131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12133 = 9'h161 == r_count_29_io_out ? io_r_353_b : _GEN_12132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12134 = 9'h162 == r_count_29_io_out ? io_r_354_b : _GEN_12133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12135 = 9'h163 == r_count_29_io_out ? io_r_355_b : _GEN_12134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12136 = 9'h164 == r_count_29_io_out ? io_r_356_b : _GEN_12135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12137 = 9'h165 == r_count_29_io_out ? io_r_357_b : _GEN_12136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12138 = 9'h166 == r_count_29_io_out ? io_r_358_b : _GEN_12137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12139 = 9'h167 == r_count_29_io_out ? io_r_359_b : _GEN_12138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12140 = 9'h168 == r_count_29_io_out ? io_r_360_b : _GEN_12139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12141 = 9'h169 == r_count_29_io_out ? io_r_361_b : _GEN_12140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12142 = 9'h16a == r_count_29_io_out ? io_r_362_b : _GEN_12141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12143 = 9'h16b == r_count_29_io_out ? io_r_363_b : _GEN_12142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12144 = 9'h16c == r_count_29_io_out ? io_r_364_b : _GEN_12143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12145 = 9'h16d == r_count_29_io_out ? io_r_365_b : _GEN_12144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12146 = 9'h16e == r_count_29_io_out ? io_r_366_b : _GEN_12145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12147 = 9'h16f == r_count_29_io_out ? io_r_367_b : _GEN_12146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12148 = 9'h170 == r_count_29_io_out ? io_r_368_b : _GEN_12147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12149 = 9'h171 == r_count_29_io_out ? io_r_369_b : _GEN_12148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12150 = 9'h172 == r_count_29_io_out ? io_r_370_b : _GEN_12149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12151 = 9'h173 == r_count_29_io_out ? io_r_371_b : _GEN_12150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12152 = 9'h174 == r_count_29_io_out ? io_r_372_b : _GEN_12151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12153 = 9'h175 == r_count_29_io_out ? io_r_373_b : _GEN_12152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12154 = 9'h176 == r_count_29_io_out ? io_r_374_b : _GEN_12153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12155 = 9'h177 == r_count_29_io_out ? io_r_375_b : _GEN_12154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12156 = 9'h178 == r_count_29_io_out ? io_r_376_b : _GEN_12155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12157 = 9'h179 == r_count_29_io_out ? io_r_377_b : _GEN_12156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12158 = 9'h17a == r_count_29_io_out ? io_r_378_b : _GEN_12157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12159 = 9'h17b == r_count_29_io_out ? io_r_379_b : _GEN_12158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12160 = 9'h17c == r_count_29_io_out ? io_r_380_b : _GEN_12159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12161 = 9'h17d == r_count_29_io_out ? io_r_381_b : _GEN_12160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12162 = 9'h17e == r_count_29_io_out ? io_r_382_b : _GEN_12161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12163 = 9'h17f == r_count_29_io_out ? io_r_383_b : _GEN_12162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12164 = 9'h180 == r_count_29_io_out ? io_r_384_b : _GEN_12163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12165 = 9'h181 == r_count_29_io_out ? io_r_385_b : _GEN_12164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12166 = 9'h182 == r_count_29_io_out ? io_r_386_b : _GEN_12165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12167 = 9'h183 == r_count_29_io_out ? io_r_387_b : _GEN_12166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12168 = 9'h184 == r_count_29_io_out ? io_r_388_b : _GEN_12167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12169 = 9'h185 == r_count_29_io_out ? io_r_389_b : _GEN_12168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12170 = 9'h186 == r_count_29_io_out ? io_r_390_b : _GEN_12169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12171 = 9'h187 == r_count_29_io_out ? io_r_391_b : _GEN_12170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12172 = 9'h188 == r_count_29_io_out ? io_r_392_b : _GEN_12171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12173 = 9'h189 == r_count_29_io_out ? io_r_393_b : _GEN_12172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12174 = 9'h18a == r_count_29_io_out ? io_r_394_b : _GEN_12173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12175 = 9'h18b == r_count_29_io_out ? io_r_395_b : _GEN_12174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12176 = 9'h18c == r_count_29_io_out ? io_r_396_b : _GEN_12175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12177 = 9'h18d == r_count_29_io_out ? io_r_397_b : _GEN_12176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12178 = 9'h18e == r_count_29_io_out ? io_r_398_b : _GEN_12177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12181 = 9'h1 == r_count_30_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12182 = 9'h2 == r_count_30_io_out ? io_r_2_b : _GEN_12181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12183 = 9'h3 == r_count_30_io_out ? io_r_3_b : _GEN_12182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12184 = 9'h4 == r_count_30_io_out ? io_r_4_b : _GEN_12183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12185 = 9'h5 == r_count_30_io_out ? io_r_5_b : _GEN_12184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12186 = 9'h6 == r_count_30_io_out ? io_r_6_b : _GEN_12185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12187 = 9'h7 == r_count_30_io_out ? io_r_7_b : _GEN_12186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12188 = 9'h8 == r_count_30_io_out ? io_r_8_b : _GEN_12187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12189 = 9'h9 == r_count_30_io_out ? io_r_9_b : _GEN_12188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12190 = 9'ha == r_count_30_io_out ? io_r_10_b : _GEN_12189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12191 = 9'hb == r_count_30_io_out ? io_r_11_b : _GEN_12190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12192 = 9'hc == r_count_30_io_out ? io_r_12_b : _GEN_12191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12193 = 9'hd == r_count_30_io_out ? io_r_13_b : _GEN_12192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12194 = 9'he == r_count_30_io_out ? io_r_14_b : _GEN_12193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12195 = 9'hf == r_count_30_io_out ? io_r_15_b : _GEN_12194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12196 = 9'h10 == r_count_30_io_out ? io_r_16_b : _GEN_12195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12197 = 9'h11 == r_count_30_io_out ? io_r_17_b : _GEN_12196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12198 = 9'h12 == r_count_30_io_out ? io_r_18_b : _GEN_12197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12199 = 9'h13 == r_count_30_io_out ? io_r_19_b : _GEN_12198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12200 = 9'h14 == r_count_30_io_out ? io_r_20_b : _GEN_12199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12201 = 9'h15 == r_count_30_io_out ? io_r_21_b : _GEN_12200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12202 = 9'h16 == r_count_30_io_out ? io_r_22_b : _GEN_12201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12203 = 9'h17 == r_count_30_io_out ? io_r_23_b : _GEN_12202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12204 = 9'h18 == r_count_30_io_out ? io_r_24_b : _GEN_12203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12205 = 9'h19 == r_count_30_io_out ? io_r_25_b : _GEN_12204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12206 = 9'h1a == r_count_30_io_out ? io_r_26_b : _GEN_12205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12207 = 9'h1b == r_count_30_io_out ? io_r_27_b : _GEN_12206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12208 = 9'h1c == r_count_30_io_out ? io_r_28_b : _GEN_12207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12209 = 9'h1d == r_count_30_io_out ? io_r_29_b : _GEN_12208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12210 = 9'h1e == r_count_30_io_out ? io_r_30_b : _GEN_12209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12211 = 9'h1f == r_count_30_io_out ? io_r_31_b : _GEN_12210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12212 = 9'h20 == r_count_30_io_out ? io_r_32_b : _GEN_12211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12213 = 9'h21 == r_count_30_io_out ? io_r_33_b : _GEN_12212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12214 = 9'h22 == r_count_30_io_out ? io_r_34_b : _GEN_12213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12215 = 9'h23 == r_count_30_io_out ? io_r_35_b : _GEN_12214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12216 = 9'h24 == r_count_30_io_out ? io_r_36_b : _GEN_12215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12217 = 9'h25 == r_count_30_io_out ? io_r_37_b : _GEN_12216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12218 = 9'h26 == r_count_30_io_out ? io_r_38_b : _GEN_12217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12219 = 9'h27 == r_count_30_io_out ? io_r_39_b : _GEN_12218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12220 = 9'h28 == r_count_30_io_out ? io_r_40_b : _GEN_12219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12221 = 9'h29 == r_count_30_io_out ? io_r_41_b : _GEN_12220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12222 = 9'h2a == r_count_30_io_out ? io_r_42_b : _GEN_12221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12223 = 9'h2b == r_count_30_io_out ? io_r_43_b : _GEN_12222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12224 = 9'h2c == r_count_30_io_out ? io_r_44_b : _GEN_12223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12225 = 9'h2d == r_count_30_io_out ? io_r_45_b : _GEN_12224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12226 = 9'h2e == r_count_30_io_out ? io_r_46_b : _GEN_12225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12227 = 9'h2f == r_count_30_io_out ? io_r_47_b : _GEN_12226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12228 = 9'h30 == r_count_30_io_out ? io_r_48_b : _GEN_12227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12229 = 9'h31 == r_count_30_io_out ? io_r_49_b : _GEN_12228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12230 = 9'h32 == r_count_30_io_out ? io_r_50_b : _GEN_12229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12231 = 9'h33 == r_count_30_io_out ? io_r_51_b : _GEN_12230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12232 = 9'h34 == r_count_30_io_out ? io_r_52_b : _GEN_12231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12233 = 9'h35 == r_count_30_io_out ? io_r_53_b : _GEN_12232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12234 = 9'h36 == r_count_30_io_out ? io_r_54_b : _GEN_12233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12235 = 9'h37 == r_count_30_io_out ? io_r_55_b : _GEN_12234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12236 = 9'h38 == r_count_30_io_out ? io_r_56_b : _GEN_12235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12237 = 9'h39 == r_count_30_io_out ? io_r_57_b : _GEN_12236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12238 = 9'h3a == r_count_30_io_out ? io_r_58_b : _GEN_12237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12239 = 9'h3b == r_count_30_io_out ? io_r_59_b : _GEN_12238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12240 = 9'h3c == r_count_30_io_out ? io_r_60_b : _GEN_12239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12241 = 9'h3d == r_count_30_io_out ? io_r_61_b : _GEN_12240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12242 = 9'h3e == r_count_30_io_out ? io_r_62_b : _GEN_12241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12243 = 9'h3f == r_count_30_io_out ? io_r_63_b : _GEN_12242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12244 = 9'h40 == r_count_30_io_out ? io_r_64_b : _GEN_12243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12245 = 9'h41 == r_count_30_io_out ? io_r_65_b : _GEN_12244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12246 = 9'h42 == r_count_30_io_out ? io_r_66_b : _GEN_12245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12247 = 9'h43 == r_count_30_io_out ? io_r_67_b : _GEN_12246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12248 = 9'h44 == r_count_30_io_out ? io_r_68_b : _GEN_12247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12249 = 9'h45 == r_count_30_io_out ? io_r_69_b : _GEN_12248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12250 = 9'h46 == r_count_30_io_out ? io_r_70_b : _GEN_12249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12251 = 9'h47 == r_count_30_io_out ? io_r_71_b : _GEN_12250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12252 = 9'h48 == r_count_30_io_out ? io_r_72_b : _GEN_12251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12253 = 9'h49 == r_count_30_io_out ? io_r_73_b : _GEN_12252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12254 = 9'h4a == r_count_30_io_out ? io_r_74_b : _GEN_12253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12255 = 9'h4b == r_count_30_io_out ? io_r_75_b : _GEN_12254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12256 = 9'h4c == r_count_30_io_out ? io_r_76_b : _GEN_12255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12257 = 9'h4d == r_count_30_io_out ? io_r_77_b : _GEN_12256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12258 = 9'h4e == r_count_30_io_out ? io_r_78_b : _GEN_12257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12259 = 9'h4f == r_count_30_io_out ? io_r_79_b : _GEN_12258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12260 = 9'h50 == r_count_30_io_out ? io_r_80_b : _GEN_12259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12261 = 9'h51 == r_count_30_io_out ? io_r_81_b : _GEN_12260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12262 = 9'h52 == r_count_30_io_out ? io_r_82_b : _GEN_12261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12263 = 9'h53 == r_count_30_io_out ? io_r_83_b : _GEN_12262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12264 = 9'h54 == r_count_30_io_out ? io_r_84_b : _GEN_12263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12265 = 9'h55 == r_count_30_io_out ? io_r_85_b : _GEN_12264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12266 = 9'h56 == r_count_30_io_out ? io_r_86_b : _GEN_12265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12267 = 9'h57 == r_count_30_io_out ? io_r_87_b : _GEN_12266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12268 = 9'h58 == r_count_30_io_out ? io_r_88_b : _GEN_12267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12269 = 9'h59 == r_count_30_io_out ? io_r_89_b : _GEN_12268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12270 = 9'h5a == r_count_30_io_out ? io_r_90_b : _GEN_12269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12271 = 9'h5b == r_count_30_io_out ? io_r_91_b : _GEN_12270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12272 = 9'h5c == r_count_30_io_out ? io_r_92_b : _GEN_12271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12273 = 9'h5d == r_count_30_io_out ? io_r_93_b : _GEN_12272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12274 = 9'h5e == r_count_30_io_out ? io_r_94_b : _GEN_12273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12275 = 9'h5f == r_count_30_io_out ? io_r_95_b : _GEN_12274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12276 = 9'h60 == r_count_30_io_out ? io_r_96_b : _GEN_12275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12277 = 9'h61 == r_count_30_io_out ? io_r_97_b : _GEN_12276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12278 = 9'h62 == r_count_30_io_out ? io_r_98_b : _GEN_12277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12279 = 9'h63 == r_count_30_io_out ? io_r_99_b : _GEN_12278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12280 = 9'h64 == r_count_30_io_out ? io_r_100_b : _GEN_12279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12281 = 9'h65 == r_count_30_io_out ? io_r_101_b : _GEN_12280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12282 = 9'h66 == r_count_30_io_out ? io_r_102_b : _GEN_12281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12283 = 9'h67 == r_count_30_io_out ? io_r_103_b : _GEN_12282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12284 = 9'h68 == r_count_30_io_out ? io_r_104_b : _GEN_12283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12285 = 9'h69 == r_count_30_io_out ? io_r_105_b : _GEN_12284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12286 = 9'h6a == r_count_30_io_out ? io_r_106_b : _GEN_12285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12287 = 9'h6b == r_count_30_io_out ? io_r_107_b : _GEN_12286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12288 = 9'h6c == r_count_30_io_out ? io_r_108_b : _GEN_12287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12289 = 9'h6d == r_count_30_io_out ? io_r_109_b : _GEN_12288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12290 = 9'h6e == r_count_30_io_out ? io_r_110_b : _GEN_12289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12291 = 9'h6f == r_count_30_io_out ? io_r_111_b : _GEN_12290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12292 = 9'h70 == r_count_30_io_out ? io_r_112_b : _GEN_12291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12293 = 9'h71 == r_count_30_io_out ? io_r_113_b : _GEN_12292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12294 = 9'h72 == r_count_30_io_out ? io_r_114_b : _GEN_12293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12295 = 9'h73 == r_count_30_io_out ? io_r_115_b : _GEN_12294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12296 = 9'h74 == r_count_30_io_out ? io_r_116_b : _GEN_12295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12297 = 9'h75 == r_count_30_io_out ? io_r_117_b : _GEN_12296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12298 = 9'h76 == r_count_30_io_out ? io_r_118_b : _GEN_12297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12299 = 9'h77 == r_count_30_io_out ? io_r_119_b : _GEN_12298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12300 = 9'h78 == r_count_30_io_out ? io_r_120_b : _GEN_12299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12301 = 9'h79 == r_count_30_io_out ? io_r_121_b : _GEN_12300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12302 = 9'h7a == r_count_30_io_out ? io_r_122_b : _GEN_12301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12303 = 9'h7b == r_count_30_io_out ? io_r_123_b : _GEN_12302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12304 = 9'h7c == r_count_30_io_out ? io_r_124_b : _GEN_12303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12305 = 9'h7d == r_count_30_io_out ? io_r_125_b : _GEN_12304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12306 = 9'h7e == r_count_30_io_out ? io_r_126_b : _GEN_12305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12307 = 9'h7f == r_count_30_io_out ? io_r_127_b : _GEN_12306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12308 = 9'h80 == r_count_30_io_out ? io_r_128_b : _GEN_12307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12309 = 9'h81 == r_count_30_io_out ? io_r_129_b : _GEN_12308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12310 = 9'h82 == r_count_30_io_out ? io_r_130_b : _GEN_12309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12311 = 9'h83 == r_count_30_io_out ? io_r_131_b : _GEN_12310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12312 = 9'h84 == r_count_30_io_out ? io_r_132_b : _GEN_12311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12313 = 9'h85 == r_count_30_io_out ? io_r_133_b : _GEN_12312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12314 = 9'h86 == r_count_30_io_out ? io_r_134_b : _GEN_12313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12315 = 9'h87 == r_count_30_io_out ? io_r_135_b : _GEN_12314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12316 = 9'h88 == r_count_30_io_out ? io_r_136_b : _GEN_12315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12317 = 9'h89 == r_count_30_io_out ? io_r_137_b : _GEN_12316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12318 = 9'h8a == r_count_30_io_out ? io_r_138_b : _GEN_12317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12319 = 9'h8b == r_count_30_io_out ? io_r_139_b : _GEN_12318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12320 = 9'h8c == r_count_30_io_out ? io_r_140_b : _GEN_12319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12321 = 9'h8d == r_count_30_io_out ? io_r_141_b : _GEN_12320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12322 = 9'h8e == r_count_30_io_out ? io_r_142_b : _GEN_12321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12323 = 9'h8f == r_count_30_io_out ? io_r_143_b : _GEN_12322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12324 = 9'h90 == r_count_30_io_out ? io_r_144_b : _GEN_12323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12325 = 9'h91 == r_count_30_io_out ? io_r_145_b : _GEN_12324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12326 = 9'h92 == r_count_30_io_out ? io_r_146_b : _GEN_12325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12327 = 9'h93 == r_count_30_io_out ? io_r_147_b : _GEN_12326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12328 = 9'h94 == r_count_30_io_out ? io_r_148_b : _GEN_12327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12329 = 9'h95 == r_count_30_io_out ? io_r_149_b : _GEN_12328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12330 = 9'h96 == r_count_30_io_out ? io_r_150_b : _GEN_12329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12331 = 9'h97 == r_count_30_io_out ? io_r_151_b : _GEN_12330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12332 = 9'h98 == r_count_30_io_out ? io_r_152_b : _GEN_12331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12333 = 9'h99 == r_count_30_io_out ? io_r_153_b : _GEN_12332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12334 = 9'h9a == r_count_30_io_out ? io_r_154_b : _GEN_12333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12335 = 9'h9b == r_count_30_io_out ? io_r_155_b : _GEN_12334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12336 = 9'h9c == r_count_30_io_out ? io_r_156_b : _GEN_12335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12337 = 9'h9d == r_count_30_io_out ? io_r_157_b : _GEN_12336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12338 = 9'h9e == r_count_30_io_out ? io_r_158_b : _GEN_12337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12339 = 9'h9f == r_count_30_io_out ? io_r_159_b : _GEN_12338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12340 = 9'ha0 == r_count_30_io_out ? io_r_160_b : _GEN_12339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12341 = 9'ha1 == r_count_30_io_out ? io_r_161_b : _GEN_12340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12342 = 9'ha2 == r_count_30_io_out ? io_r_162_b : _GEN_12341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12343 = 9'ha3 == r_count_30_io_out ? io_r_163_b : _GEN_12342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12344 = 9'ha4 == r_count_30_io_out ? io_r_164_b : _GEN_12343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12345 = 9'ha5 == r_count_30_io_out ? io_r_165_b : _GEN_12344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12346 = 9'ha6 == r_count_30_io_out ? io_r_166_b : _GEN_12345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12347 = 9'ha7 == r_count_30_io_out ? io_r_167_b : _GEN_12346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12348 = 9'ha8 == r_count_30_io_out ? io_r_168_b : _GEN_12347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12349 = 9'ha9 == r_count_30_io_out ? io_r_169_b : _GEN_12348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12350 = 9'haa == r_count_30_io_out ? io_r_170_b : _GEN_12349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12351 = 9'hab == r_count_30_io_out ? io_r_171_b : _GEN_12350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12352 = 9'hac == r_count_30_io_out ? io_r_172_b : _GEN_12351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12353 = 9'had == r_count_30_io_out ? io_r_173_b : _GEN_12352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12354 = 9'hae == r_count_30_io_out ? io_r_174_b : _GEN_12353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12355 = 9'haf == r_count_30_io_out ? io_r_175_b : _GEN_12354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12356 = 9'hb0 == r_count_30_io_out ? io_r_176_b : _GEN_12355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12357 = 9'hb1 == r_count_30_io_out ? io_r_177_b : _GEN_12356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12358 = 9'hb2 == r_count_30_io_out ? io_r_178_b : _GEN_12357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12359 = 9'hb3 == r_count_30_io_out ? io_r_179_b : _GEN_12358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12360 = 9'hb4 == r_count_30_io_out ? io_r_180_b : _GEN_12359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12361 = 9'hb5 == r_count_30_io_out ? io_r_181_b : _GEN_12360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12362 = 9'hb6 == r_count_30_io_out ? io_r_182_b : _GEN_12361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12363 = 9'hb7 == r_count_30_io_out ? io_r_183_b : _GEN_12362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12364 = 9'hb8 == r_count_30_io_out ? io_r_184_b : _GEN_12363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12365 = 9'hb9 == r_count_30_io_out ? io_r_185_b : _GEN_12364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12366 = 9'hba == r_count_30_io_out ? io_r_186_b : _GEN_12365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12367 = 9'hbb == r_count_30_io_out ? io_r_187_b : _GEN_12366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12368 = 9'hbc == r_count_30_io_out ? io_r_188_b : _GEN_12367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12369 = 9'hbd == r_count_30_io_out ? io_r_189_b : _GEN_12368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12370 = 9'hbe == r_count_30_io_out ? io_r_190_b : _GEN_12369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12371 = 9'hbf == r_count_30_io_out ? io_r_191_b : _GEN_12370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12372 = 9'hc0 == r_count_30_io_out ? io_r_192_b : _GEN_12371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12373 = 9'hc1 == r_count_30_io_out ? io_r_193_b : _GEN_12372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12374 = 9'hc2 == r_count_30_io_out ? io_r_194_b : _GEN_12373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12375 = 9'hc3 == r_count_30_io_out ? io_r_195_b : _GEN_12374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12376 = 9'hc4 == r_count_30_io_out ? io_r_196_b : _GEN_12375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12377 = 9'hc5 == r_count_30_io_out ? io_r_197_b : _GEN_12376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12378 = 9'hc6 == r_count_30_io_out ? io_r_198_b : _GEN_12377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12379 = 9'hc7 == r_count_30_io_out ? io_r_199_b : _GEN_12378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12380 = 9'hc8 == r_count_30_io_out ? io_r_200_b : _GEN_12379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12381 = 9'hc9 == r_count_30_io_out ? io_r_201_b : _GEN_12380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12382 = 9'hca == r_count_30_io_out ? io_r_202_b : _GEN_12381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12383 = 9'hcb == r_count_30_io_out ? io_r_203_b : _GEN_12382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12384 = 9'hcc == r_count_30_io_out ? io_r_204_b : _GEN_12383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12385 = 9'hcd == r_count_30_io_out ? io_r_205_b : _GEN_12384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12386 = 9'hce == r_count_30_io_out ? io_r_206_b : _GEN_12385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12387 = 9'hcf == r_count_30_io_out ? io_r_207_b : _GEN_12386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12388 = 9'hd0 == r_count_30_io_out ? io_r_208_b : _GEN_12387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12389 = 9'hd1 == r_count_30_io_out ? io_r_209_b : _GEN_12388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12390 = 9'hd2 == r_count_30_io_out ? io_r_210_b : _GEN_12389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12391 = 9'hd3 == r_count_30_io_out ? io_r_211_b : _GEN_12390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12392 = 9'hd4 == r_count_30_io_out ? io_r_212_b : _GEN_12391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12393 = 9'hd5 == r_count_30_io_out ? io_r_213_b : _GEN_12392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12394 = 9'hd6 == r_count_30_io_out ? io_r_214_b : _GEN_12393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12395 = 9'hd7 == r_count_30_io_out ? io_r_215_b : _GEN_12394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12396 = 9'hd8 == r_count_30_io_out ? io_r_216_b : _GEN_12395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12397 = 9'hd9 == r_count_30_io_out ? io_r_217_b : _GEN_12396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12398 = 9'hda == r_count_30_io_out ? io_r_218_b : _GEN_12397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12399 = 9'hdb == r_count_30_io_out ? io_r_219_b : _GEN_12398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12400 = 9'hdc == r_count_30_io_out ? io_r_220_b : _GEN_12399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12401 = 9'hdd == r_count_30_io_out ? io_r_221_b : _GEN_12400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12402 = 9'hde == r_count_30_io_out ? io_r_222_b : _GEN_12401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12403 = 9'hdf == r_count_30_io_out ? io_r_223_b : _GEN_12402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12404 = 9'he0 == r_count_30_io_out ? io_r_224_b : _GEN_12403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12405 = 9'he1 == r_count_30_io_out ? io_r_225_b : _GEN_12404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12406 = 9'he2 == r_count_30_io_out ? io_r_226_b : _GEN_12405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12407 = 9'he3 == r_count_30_io_out ? io_r_227_b : _GEN_12406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12408 = 9'he4 == r_count_30_io_out ? io_r_228_b : _GEN_12407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12409 = 9'he5 == r_count_30_io_out ? io_r_229_b : _GEN_12408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12410 = 9'he6 == r_count_30_io_out ? io_r_230_b : _GEN_12409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12411 = 9'he7 == r_count_30_io_out ? io_r_231_b : _GEN_12410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12412 = 9'he8 == r_count_30_io_out ? io_r_232_b : _GEN_12411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12413 = 9'he9 == r_count_30_io_out ? io_r_233_b : _GEN_12412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12414 = 9'hea == r_count_30_io_out ? io_r_234_b : _GEN_12413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12415 = 9'heb == r_count_30_io_out ? io_r_235_b : _GEN_12414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12416 = 9'hec == r_count_30_io_out ? io_r_236_b : _GEN_12415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12417 = 9'hed == r_count_30_io_out ? io_r_237_b : _GEN_12416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12418 = 9'hee == r_count_30_io_out ? io_r_238_b : _GEN_12417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12419 = 9'hef == r_count_30_io_out ? io_r_239_b : _GEN_12418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12420 = 9'hf0 == r_count_30_io_out ? io_r_240_b : _GEN_12419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12421 = 9'hf1 == r_count_30_io_out ? io_r_241_b : _GEN_12420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12422 = 9'hf2 == r_count_30_io_out ? io_r_242_b : _GEN_12421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12423 = 9'hf3 == r_count_30_io_out ? io_r_243_b : _GEN_12422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12424 = 9'hf4 == r_count_30_io_out ? io_r_244_b : _GEN_12423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12425 = 9'hf5 == r_count_30_io_out ? io_r_245_b : _GEN_12424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12426 = 9'hf6 == r_count_30_io_out ? io_r_246_b : _GEN_12425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12427 = 9'hf7 == r_count_30_io_out ? io_r_247_b : _GEN_12426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12428 = 9'hf8 == r_count_30_io_out ? io_r_248_b : _GEN_12427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12429 = 9'hf9 == r_count_30_io_out ? io_r_249_b : _GEN_12428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12430 = 9'hfa == r_count_30_io_out ? io_r_250_b : _GEN_12429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12431 = 9'hfb == r_count_30_io_out ? io_r_251_b : _GEN_12430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12432 = 9'hfc == r_count_30_io_out ? io_r_252_b : _GEN_12431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12433 = 9'hfd == r_count_30_io_out ? io_r_253_b : _GEN_12432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12434 = 9'hfe == r_count_30_io_out ? io_r_254_b : _GEN_12433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12435 = 9'hff == r_count_30_io_out ? io_r_255_b : _GEN_12434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12436 = 9'h100 == r_count_30_io_out ? io_r_256_b : _GEN_12435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12437 = 9'h101 == r_count_30_io_out ? io_r_257_b : _GEN_12436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12438 = 9'h102 == r_count_30_io_out ? io_r_258_b : _GEN_12437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12439 = 9'h103 == r_count_30_io_out ? io_r_259_b : _GEN_12438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12440 = 9'h104 == r_count_30_io_out ? io_r_260_b : _GEN_12439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12441 = 9'h105 == r_count_30_io_out ? io_r_261_b : _GEN_12440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12442 = 9'h106 == r_count_30_io_out ? io_r_262_b : _GEN_12441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12443 = 9'h107 == r_count_30_io_out ? io_r_263_b : _GEN_12442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12444 = 9'h108 == r_count_30_io_out ? io_r_264_b : _GEN_12443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12445 = 9'h109 == r_count_30_io_out ? io_r_265_b : _GEN_12444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12446 = 9'h10a == r_count_30_io_out ? io_r_266_b : _GEN_12445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12447 = 9'h10b == r_count_30_io_out ? io_r_267_b : _GEN_12446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12448 = 9'h10c == r_count_30_io_out ? io_r_268_b : _GEN_12447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12449 = 9'h10d == r_count_30_io_out ? io_r_269_b : _GEN_12448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12450 = 9'h10e == r_count_30_io_out ? io_r_270_b : _GEN_12449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12451 = 9'h10f == r_count_30_io_out ? io_r_271_b : _GEN_12450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12452 = 9'h110 == r_count_30_io_out ? io_r_272_b : _GEN_12451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12453 = 9'h111 == r_count_30_io_out ? io_r_273_b : _GEN_12452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12454 = 9'h112 == r_count_30_io_out ? io_r_274_b : _GEN_12453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12455 = 9'h113 == r_count_30_io_out ? io_r_275_b : _GEN_12454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12456 = 9'h114 == r_count_30_io_out ? io_r_276_b : _GEN_12455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12457 = 9'h115 == r_count_30_io_out ? io_r_277_b : _GEN_12456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12458 = 9'h116 == r_count_30_io_out ? io_r_278_b : _GEN_12457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12459 = 9'h117 == r_count_30_io_out ? io_r_279_b : _GEN_12458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12460 = 9'h118 == r_count_30_io_out ? io_r_280_b : _GEN_12459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12461 = 9'h119 == r_count_30_io_out ? io_r_281_b : _GEN_12460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12462 = 9'h11a == r_count_30_io_out ? io_r_282_b : _GEN_12461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12463 = 9'h11b == r_count_30_io_out ? io_r_283_b : _GEN_12462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12464 = 9'h11c == r_count_30_io_out ? io_r_284_b : _GEN_12463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12465 = 9'h11d == r_count_30_io_out ? io_r_285_b : _GEN_12464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12466 = 9'h11e == r_count_30_io_out ? io_r_286_b : _GEN_12465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12467 = 9'h11f == r_count_30_io_out ? io_r_287_b : _GEN_12466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12468 = 9'h120 == r_count_30_io_out ? io_r_288_b : _GEN_12467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12469 = 9'h121 == r_count_30_io_out ? io_r_289_b : _GEN_12468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12470 = 9'h122 == r_count_30_io_out ? io_r_290_b : _GEN_12469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12471 = 9'h123 == r_count_30_io_out ? io_r_291_b : _GEN_12470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12472 = 9'h124 == r_count_30_io_out ? io_r_292_b : _GEN_12471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12473 = 9'h125 == r_count_30_io_out ? io_r_293_b : _GEN_12472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12474 = 9'h126 == r_count_30_io_out ? io_r_294_b : _GEN_12473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12475 = 9'h127 == r_count_30_io_out ? io_r_295_b : _GEN_12474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12476 = 9'h128 == r_count_30_io_out ? io_r_296_b : _GEN_12475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12477 = 9'h129 == r_count_30_io_out ? io_r_297_b : _GEN_12476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12478 = 9'h12a == r_count_30_io_out ? io_r_298_b : _GEN_12477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12479 = 9'h12b == r_count_30_io_out ? io_r_299_b : _GEN_12478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12480 = 9'h12c == r_count_30_io_out ? io_r_300_b : _GEN_12479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12481 = 9'h12d == r_count_30_io_out ? io_r_301_b : _GEN_12480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12482 = 9'h12e == r_count_30_io_out ? io_r_302_b : _GEN_12481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12483 = 9'h12f == r_count_30_io_out ? io_r_303_b : _GEN_12482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12484 = 9'h130 == r_count_30_io_out ? io_r_304_b : _GEN_12483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12485 = 9'h131 == r_count_30_io_out ? io_r_305_b : _GEN_12484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12486 = 9'h132 == r_count_30_io_out ? io_r_306_b : _GEN_12485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12487 = 9'h133 == r_count_30_io_out ? io_r_307_b : _GEN_12486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12488 = 9'h134 == r_count_30_io_out ? io_r_308_b : _GEN_12487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12489 = 9'h135 == r_count_30_io_out ? io_r_309_b : _GEN_12488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12490 = 9'h136 == r_count_30_io_out ? io_r_310_b : _GEN_12489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12491 = 9'h137 == r_count_30_io_out ? io_r_311_b : _GEN_12490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12492 = 9'h138 == r_count_30_io_out ? io_r_312_b : _GEN_12491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12493 = 9'h139 == r_count_30_io_out ? io_r_313_b : _GEN_12492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12494 = 9'h13a == r_count_30_io_out ? io_r_314_b : _GEN_12493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12495 = 9'h13b == r_count_30_io_out ? io_r_315_b : _GEN_12494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12496 = 9'h13c == r_count_30_io_out ? io_r_316_b : _GEN_12495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12497 = 9'h13d == r_count_30_io_out ? io_r_317_b : _GEN_12496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12498 = 9'h13e == r_count_30_io_out ? io_r_318_b : _GEN_12497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12499 = 9'h13f == r_count_30_io_out ? io_r_319_b : _GEN_12498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12500 = 9'h140 == r_count_30_io_out ? io_r_320_b : _GEN_12499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12501 = 9'h141 == r_count_30_io_out ? io_r_321_b : _GEN_12500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12502 = 9'h142 == r_count_30_io_out ? io_r_322_b : _GEN_12501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12503 = 9'h143 == r_count_30_io_out ? io_r_323_b : _GEN_12502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12504 = 9'h144 == r_count_30_io_out ? io_r_324_b : _GEN_12503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12505 = 9'h145 == r_count_30_io_out ? io_r_325_b : _GEN_12504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12506 = 9'h146 == r_count_30_io_out ? io_r_326_b : _GEN_12505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12507 = 9'h147 == r_count_30_io_out ? io_r_327_b : _GEN_12506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12508 = 9'h148 == r_count_30_io_out ? io_r_328_b : _GEN_12507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12509 = 9'h149 == r_count_30_io_out ? io_r_329_b : _GEN_12508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12510 = 9'h14a == r_count_30_io_out ? io_r_330_b : _GEN_12509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12511 = 9'h14b == r_count_30_io_out ? io_r_331_b : _GEN_12510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12512 = 9'h14c == r_count_30_io_out ? io_r_332_b : _GEN_12511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12513 = 9'h14d == r_count_30_io_out ? io_r_333_b : _GEN_12512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12514 = 9'h14e == r_count_30_io_out ? io_r_334_b : _GEN_12513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12515 = 9'h14f == r_count_30_io_out ? io_r_335_b : _GEN_12514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12516 = 9'h150 == r_count_30_io_out ? io_r_336_b : _GEN_12515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12517 = 9'h151 == r_count_30_io_out ? io_r_337_b : _GEN_12516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12518 = 9'h152 == r_count_30_io_out ? io_r_338_b : _GEN_12517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12519 = 9'h153 == r_count_30_io_out ? io_r_339_b : _GEN_12518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12520 = 9'h154 == r_count_30_io_out ? io_r_340_b : _GEN_12519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12521 = 9'h155 == r_count_30_io_out ? io_r_341_b : _GEN_12520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12522 = 9'h156 == r_count_30_io_out ? io_r_342_b : _GEN_12521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12523 = 9'h157 == r_count_30_io_out ? io_r_343_b : _GEN_12522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12524 = 9'h158 == r_count_30_io_out ? io_r_344_b : _GEN_12523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12525 = 9'h159 == r_count_30_io_out ? io_r_345_b : _GEN_12524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12526 = 9'h15a == r_count_30_io_out ? io_r_346_b : _GEN_12525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12527 = 9'h15b == r_count_30_io_out ? io_r_347_b : _GEN_12526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12528 = 9'h15c == r_count_30_io_out ? io_r_348_b : _GEN_12527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12529 = 9'h15d == r_count_30_io_out ? io_r_349_b : _GEN_12528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12530 = 9'h15e == r_count_30_io_out ? io_r_350_b : _GEN_12529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12531 = 9'h15f == r_count_30_io_out ? io_r_351_b : _GEN_12530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12532 = 9'h160 == r_count_30_io_out ? io_r_352_b : _GEN_12531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12533 = 9'h161 == r_count_30_io_out ? io_r_353_b : _GEN_12532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12534 = 9'h162 == r_count_30_io_out ? io_r_354_b : _GEN_12533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12535 = 9'h163 == r_count_30_io_out ? io_r_355_b : _GEN_12534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12536 = 9'h164 == r_count_30_io_out ? io_r_356_b : _GEN_12535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12537 = 9'h165 == r_count_30_io_out ? io_r_357_b : _GEN_12536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12538 = 9'h166 == r_count_30_io_out ? io_r_358_b : _GEN_12537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12539 = 9'h167 == r_count_30_io_out ? io_r_359_b : _GEN_12538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12540 = 9'h168 == r_count_30_io_out ? io_r_360_b : _GEN_12539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12541 = 9'h169 == r_count_30_io_out ? io_r_361_b : _GEN_12540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12542 = 9'h16a == r_count_30_io_out ? io_r_362_b : _GEN_12541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12543 = 9'h16b == r_count_30_io_out ? io_r_363_b : _GEN_12542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12544 = 9'h16c == r_count_30_io_out ? io_r_364_b : _GEN_12543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12545 = 9'h16d == r_count_30_io_out ? io_r_365_b : _GEN_12544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12546 = 9'h16e == r_count_30_io_out ? io_r_366_b : _GEN_12545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12547 = 9'h16f == r_count_30_io_out ? io_r_367_b : _GEN_12546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12548 = 9'h170 == r_count_30_io_out ? io_r_368_b : _GEN_12547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12549 = 9'h171 == r_count_30_io_out ? io_r_369_b : _GEN_12548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12550 = 9'h172 == r_count_30_io_out ? io_r_370_b : _GEN_12549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12551 = 9'h173 == r_count_30_io_out ? io_r_371_b : _GEN_12550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12552 = 9'h174 == r_count_30_io_out ? io_r_372_b : _GEN_12551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12553 = 9'h175 == r_count_30_io_out ? io_r_373_b : _GEN_12552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12554 = 9'h176 == r_count_30_io_out ? io_r_374_b : _GEN_12553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12555 = 9'h177 == r_count_30_io_out ? io_r_375_b : _GEN_12554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12556 = 9'h178 == r_count_30_io_out ? io_r_376_b : _GEN_12555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12557 = 9'h179 == r_count_30_io_out ? io_r_377_b : _GEN_12556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12558 = 9'h17a == r_count_30_io_out ? io_r_378_b : _GEN_12557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12559 = 9'h17b == r_count_30_io_out ? io_r_379_b : _GEN_12558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12560 = 9'h17c == r_count_30_io_out ? io_r_380_b : _GEN_12559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12561 = 9'h17d == r_count_30_io_out ? io_r_381_b : _GEN_12560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12562 = 9'h17e == r_count_30_io_out ? io_r_382_b : _GEN_12561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12563 = 9'h17f == r_count_30_io_out ? io_r_383_b : _GEN_12562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12564 = 9'h180 == r_count_30_io_out ? io_r_384_b : _GEN_12563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12565 = 9'h181 == r_count_30_io_out ? io_r_385_b : _GEN_12564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12566 = 9'h182 == r_count_30_io_out ? io_r_386_b : _GEN_12565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12567 = 9'h183 == r_count_30_io_out ? io_r_387_b : _GEN_12566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12568 = 9'h184 == r_count_30_io_out ? io_r_388_b : _GEN_12567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12569 = 9'h185 == r_count_30_io_out ? io_r_389_b : _GEN_12568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12570 = 9'h186 == r_count_30_io_out ? io_r_390_b : _GEN_12569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12571 = 9'h187 == r_count_30_io_out ? io_r_391_b : _GEN_12570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12572 = 9'h188 == r_count_30_io_out ? io_r_392_b : _GEN_12571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12573 = 9'h189 == r_count_30_io_out ? io_r_393_b : _GEN_12572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12574 = 9'h18a == r_count_30_io_out ? io_r_394_b : _GEN_12573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12575 = 9'h18b == r_count_30_io_out ? io_r_395_b : _GEN_12574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12576 = 9'h18c == r_count_30_io_out ? io_r_396_b : _GEN_12575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12577 = 9'h18d == r_count_30_io_out ? io_r_397_b : _GEN_12576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12578 = 9'h18e == r_count_30_io_out ? io_r_398_b : _GEN_12577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12581 = 9'h1 == r_count_31_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12582 = 9'h2 == r_count_31_io_out ? io_r_2_b : _GEN_12581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12583 = 9'h3 == r_count_31_io_out ? io_r_3_b : _GEN_12582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12584 = 9'h4 == r_count_31_io_out ? io_r_4_b : _GEN_12583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12585 = 9'h5 == r_count_31_io_out ? io_r_5_b : _GEN_12584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12586 = 9'h6 == r_count_31_io_out ? io_r_6_b : _GEN_12585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12587 = 9'h7 == r_count_31_io_out ? io_r_7_b : _GEN_12586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12588 = 9'h8 == r_count_31_io_out ? io_r_8_b : _GEN_12587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12589 = 9'h9 == r_count_31_io_out ? io_r_9_b : _GEN_12588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12590 = 9'ha == r_count_31_io_out ? io_r_10_b : _GEN_12589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12591 = 9'hb == r_count_31_io_out ? io_r_11_b : _GEN_12590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12592 = 9'hc == r_count_31_io_out ? io_r_12_b : _GEN_12591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12593 = 9'hd == r_count_31_io_out ? io_r_13_b : _GEN_12592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12594 = 9'he == r_count_31_io_out ? io_r_14_b : _GEN_12593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12595 = 9'hf == r_count_31_io_out ? io_r_15_b : _GEN_12594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12596 = 9'h10 == r_count_31_io_out ? io_r_16_b : _GEN_12595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12597 = 9'h11 == r_count_31_io_out ? io_r_17_b : _GEN_12596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12598 = 9'h12 == r_count_31_io_out ? io_r_18_b : _GEN_12597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12599 = 9'h13 == r_count_31_io_out ? io_r_19_b : _GEN_12598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12600 = 9'h14 == r_count_31_io_out ? io_r_20_b : _GEN_12599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12601 = 9'h15 == r_count_31_io_out ? io_r_21_b : _GEN_12600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12602 = 9'h16 == r_count_31_io_out ? io_r_22_b : _GEN_12601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12603 = 9'h17 == r_count_31_io_out ? io_r_23_b : _GEN_12602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12604 = 9'h18 == r_count_31_io_out ? io_r_24_b : _GEN_12603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12605 = 9'h19 == r_count_31_io_out ? io_r_25_b : _GEN_12604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12606 = 9'h1a == r_count_31_io_out ? io_r_26_b : _GEN_12605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12607 = 9'h1b == r_count_31_io_out ? io_r_27_b : _GEN_12606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12608 = 9'h1c == r_count_31_io_out ? io_r_28_b : _GEN_12607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12609 = 9'h1d == r_count_31_io_out ? io_r_29_b : _GEN_12608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12610 = 9'h1e == r_count_31_io_out ? io_r_30_b : _GEN_12609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12611 = 9'h1f == r_count_31_io_out ? io_r_31_b : _GEN_12610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12612 = 9'h20 == r_count_31_io_out ? io_r_32_b : _GEN_12611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12613 = 9'h21 == r_count_31_io_out ? io_r_33_b : _GEN_12612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12614 = 9'h22 == r_count_31_io_out ? io_r_34_b : _GEN_12613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12615 = 9'h23 == r_count_31_io_out ? io_r_35_b : _GEN_12614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12616 = 9'h24 == r_count_31_io_out ? io_r_36_b : _GEN_12615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12617 = 9'h25 == r_count_31_io_out ? io_r_37_b : _GEN_12616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12618 = 9'h26 == r_count_31_io_out ? io_r_38_b : _GEN_12617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12619 = 9'h27 == r_count_31_io_out ? io_r_39_b : _GEN_12618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12620 = 9'h28 == r_count_31_io_out ? io_r_40_b : _GEN_12619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12621 = 9'h29 == r_count_31_io_out ? io_r_41_b : _GEN_12620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12622 = 9'h2a == r_count_31_io_out ? io_r_42_b : _GEN_12621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12623 = 9'h2b == r_count_31_io_out ? io_r_43_b : _GEN_12622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12624 = 9'h2c == r_count_31_io_out ? io_r_44_b : _GEN_12623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12625 = 9'h2d == r_count_31_io_out ? io_r_45_b : _GEN_12624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12626 = 9'h2e == r_count_31_io_out ? io_r_46_b : _GEN_12625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12627 = 9'h2f == r_count_31_io_out ? io_r_47_b : _GEN_12626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12628 = 9'h30 == r_count_31_io_out ? io_r_48_b : _GEN_12627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12629 = 9'h31 == r_count_31_io_out ? io_r_49_b : _GEN_12628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12630 = 9'h32 == r_count_31_io_out ? io_r_50_b : _GEN_12629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12631 = 9'h33 == r_count_31_io_out ? io_r_51_b : _GEN_12630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12632 = 9'h34 == r_count_31_io_out ? io_r_52_b : _GEN_12631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12633 = 9'h35 == r_count_31_io_out ? io_r_53_b : _GEN_12632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12634 = 9'h36 == r_count_31_io_out ? io_r_54_b : _GEN_12633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12635 = 9'h37 == r_count_31_io_out ? io_r_55_b : _GEN_12634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12636 = 9'h38 == r_count_31_io_out ? io_r_56_b : _GEN_12635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12637 = 9'h39 == r_count_31_io_out ? io_r_57_b : _GEN_12636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12638 = 9'h3a == r_count_31_io_out ? io_r_58_b : _GEN_12637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12639 = 9'h3b == r_count_31_io_out ? io_r_59_b : _GEN_12638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12640 = 9'h3c == r_count_31_io_out ? io_r_60_b : _GEN_12639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12641 = 9'h3d == r_count_31_io_out ? io_r_61_b : _GEN_12640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12642 = 9'h3e == r_count_31_io_out ? io_r_62_b : _GEN_12641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12643 = 9'h3f == r_count_31_io_out ? io_r_63_b : _GEN_12642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12644 = 9'h40 == r_count_31_io_out ? io_r_64_b : _GEN_12643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12645 = 9'h41 == r_count_31_io_out ? io_r_65_b : _GEN_12644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12646 = 9'h42 == r_count_31_io_out ? io_r_66_b : _GEN_12645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12647 = 9'h43 == r_count_31_io_out ? io_r_67_b : _GEN_12646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12648 = 9'h44 == r_count_31_io_out ? io_r_68_b : _GEN_12647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12649 = 9'h45 == r_count_31_io_out ? io_r_69_b : _GEN_12648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12650 = 9'h46 == r_count_31_io_out ? io_r_70_b : _GEN_12649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12651 = 9'h47 == r_count_31_io_out ? io_r_71_b : _GEN_12650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12652 = 9'h48 == r_count_31_io_out ? io_r_72_b : _GEN_12651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12653 = 9'h49 == r_count_31_io_out ? io_r_73_b : _GEN_12652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12654 = 9'h4a == r_count_31_io_out ? io_r_74_b : _GEN_12653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12655 = 9'h4b == r_count_31_io_out ? io_r_75_b : _GEN_12654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12656 = 9'h4c == r_count_31_io_out ? io_r_76_b : _GEN_12655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12657 = 9'h4d == r_count_31_io_out ? io_r_77_b : _GEN_12656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12658 = 9'h4e == r_count_31_io_out ? io_r_78_b : _GEN_12657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12659 = 9'h4f == r_count_31_io_out ? io_r_79_b : _GEN_12658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12660 = 9'h50 == r_count_31_io_out ? io_r_80_b : _GEN_12659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12661 = 9'h51 == r_count_31_io_out ? io_r_81_b : _GEN_12660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12662 = 9'h52 == r_count_31_io_out ? io_r_82_b : _GEN_12661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12663 = 9'h53 == r_count_31_io_out ? io_r_83_b : _GEN_12662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12664 = 9'h54 == r_count_31_io_out ? io_r_84_b : _GEN_12663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12665 = 9'h55 == r_count_31_io_out ? io_r_85_b : _GEN_12664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12666 = 9'h56 == r_count_31_io_out ? io_r_86_b : _GEN_12665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12667 = 9'h57 == r_count_31_io_out ? io_r_87_b : _GEN_12666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12668 = 9'h58 == r_count_31_io_out ? io_r_88_b : _GEN_12667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12669 = 9'h59 == r_count_31_io_out ? io_r_89_b : _GEN_12668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12670 = 9'h5a == r_count_31_io_out ? io_r_90_b : _GEN_12669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12671 = 9'h5b == r_count_31_io_out ? io_r_91_b : _GEN_12670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12672 = 9'h5c == r_count_31_io_out ? io_r_92_b : _GEN_12671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12673 = 9'h5d == r_count_31_io_out ? io_r_93_b : _GEN_12672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12674 = 9'h5e == r_count_31_io_out ? io_r_94_b : _GEN_12673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12675 = 9'h5f == r_count_31_io_out ? io_r_95_b : _GEN_12674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12676 = 9'h60 == r_count_31_io_out ? io_r_96_b : _GEN_12675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12677 = 9'h61 == r_count_31_io_out ? io_r_97_b : _GEN_12676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12678 = 9'h62 == r_count_31_io_out ? io_r_98_b : _GEN_12677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12679 = 9'h63 == r_count_31_io_out ? io_r_99_b : _GEN_12678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12680 = 9'h64 == r_count_31_io_out ? io_r_100_b : _GEN_12679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12681 = 9'h65 == r_count_31_io_out ? io_r_101_b : _GEN_12680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12682 = 9'h66 == r_count_31_io_out ? io_r_102_b : _GEN_12681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12683 = 9'h67 == r_count_31_io_out ? io_r_103_b : _GEN_12682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12684 = 9'h68 == r_count_31_io_out ? io_r_104_b : _GEN_12683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12685 = 9'h69 == r_count_31_io_out ? io_r_105_b : _GEN_12684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12686 = 9'h6a == r_count_31_io_out ? io_r_106_b : _GEN_12685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12687 = 9'h6b == r_count_31_io_out ? io_r_107_b : _GEN_12686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12688 = 9'h6c == r_count_31_io_out ? io_r_108_b : _GEN_12687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12689 = 9'h6d == r_count_31_io_out ? io_r_109_b : _GEN_12688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12690 = 9'h6e == r_count_31_io_out ? io_r_110_b : _GEN_12689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12691 = 9'h6f == r_count_31_io_out ? io_r_111_b : _GEN_12690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12692 = 9'h70 == r_count_31_io_out ? io_r_112_b : _GEN_12691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12693 = 9'h71 == r_count_31_io_out ? io_r_113_b : _GEN_12692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12694 = 9'h72 == r_count_31_io_out ? io_r_114_b : _GEN_12693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12695 = 9'h73 == r_count_31_io_out ? io_r_115_b : _GEN_12694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12696 = 9'h74 == r_count_31_io_out ? io_r_116_b : _GEN_12695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12697 = 9'h75 == r_count_31_io_out ? io_r_117_b : _GEN_12696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12698 = 9'h76 == r_count_31_io_out ? io_r_118_b : _GEN_12697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12699 = 9'h77 == r_count_31_io_out ? io_r_119_b : _GEN_12698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12700 = 9'h78 == r_count_31_io_out ? io_r_120_b : _GEN_12699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12701 = 9'h79 == r_count_31_io_out ? io_r_121_b : _GEN_12700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12702 = 9'h7a == r_count_31_io_out ? io_r_122_b : _GEN_12701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12703 = 9'h7b == r_count_31_io_out ? io_r_123_b : _GEN_12702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12704 = 9'h7c == r_count_31_io_out ? io_r_124_b : _GEN_12703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12705 = 9'h7d == r_count_31_io_out ? io_r_125_b : _GEN_12704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12706 = 9'h7e == r_count_31_io_out ? io_r_126_b : _GEN_12705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12707 = 9'h7f == r_count_31_io_out ? io_r_127_b : _GEN_12706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12708 = 9'h80 == r_count_31_io_out ? io_r_128_b : _GEN_12707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12709 = 9'h81 == r_count_31_io_out ? io_r_129_b : _GEN_12708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12710 = 9'h82 == r_count_31_io_out ? io_r_130_b : _GEN_12709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12711 = 9'h83 == r_count_31_io_out ? io_r_131_b : _GEN_12710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12712 = 9'h84 == r_count_31_io_out ? io_r_132_b : _GEN_12711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12713 = 9'h85 == r_count_31_io_out ? io_r_133_b : _GEN_12712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12714 = 9'h86 == r_count_31_io_out ? io_r_134_b : _GEN_12713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12715 = 9'h87 == r_count_31_io_out ? io_r_135_b : _GEN_12714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12716 = 9'h88 == r_count_31_io_out ? io_r_136_b : _GEN_12715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12717 = 9'h89 == r_count_31_io_out ? io_r_137_b : _GEN_12716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12718 = 9'h8a == r_count_31_io_out ? io_r_138_b : _GEN_12717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12719 = 9'h8b == r_count_31_io_out ? io_r_139_b : _GEN_12718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12720 = 9'h8c == r_count_31_io_out ? io_r_140_b : _GEN_12719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12721 = 9'h8d == r_count_31_io_out ? io_r_141_b : _GEN_12720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12722 = 9'h8e == r_count_31_io_out ? io_r_142_b : _GEN_12721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12723 = 9'h8f == r_count_31_io_out ? io_r_143_b : _GEN_12722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12724 = 9'h90 == r_count_31_io_out ? io_r_144_b : _GEN_12723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12725 = 9'h91 == r_count_31_io_out ? io_r_145_b : _GEN_12724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12726 = 9'h92 == r_count_31_io_out ? io_r_146_b : _GEN_12725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12727 = 9'h93 == r_count_31_io_out ? io_r_147_b : _GEN_12726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12728 = 9'h94 == r_count_31_io_out ? io_r_148_b : _GEN_12727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12729 = 9'h95 == r_count_31_io_out ? io_r_149_b : _GEN_12728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12730 = 9'h96 == r_count_31_io_out ? io_r_150_b : _GEN_12729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12731 = 9'h97 == r_count_31_io_out ? io_r_151_b : _GEN_12730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12732 = 9'h98 == r_count_31_io_out ? io_r_152_b : _GEN_12731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12733 = 9'h99 == r_count_31_io_out ? io_r_153_b : _GEN_12732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12734 = 9'h9a == r_count_31_io_out ? io_r_154_b : _GEN_12733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12735 = 9'h9b == r_count_31_io_out ? io_r_155_b : _GEN_12734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12736 = 9'h9c == r_count_31_io_out ? io_r_156_b : _GEN_12735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12737 = 9'h9d == r_count_31_io_out ? io_r_157_b : _GEN_12736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12738 = 9'h9e == r_count_31_io_out ? io_r_158_b : _GEN_12737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12739 = 9'h9f == r_count_31_io_out ? io_r_159_b : _GEN_12738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12740 = 9'ha0 == r_count_31_io_out ? io_r_160_b : _GEN_12739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12741 = 9'ha1 == r_count_31_io_out ? io_r_161_b : _GEN_12740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12742 = 9'ha2 == r_count_31_io_out ? io_r_162_b : _GEN_12741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12743 = 9'ha3 == r_count_31_io_out ? io_r_163_b : _GEN_12742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12744 = 9'ha4 == r_count_31_io_out ? io_r_164_b : _GEN_12743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12745 = 9'ha5 == r_count_31_io_out ? io_r_165_b : _GEN_12744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12746 = 9'ha6 == r_count_31_io_out ? io_r_166_b : _GEN_12745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12747 = 9'ha7 == r_count_31_io_out ? io_r_167_b : _GEN_12746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12748 = 9'ha8 == r_count_31_io_out ? io_r_168_b : _GEN_12747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12749 = 9'ha9 == r_count_31_io_out ? io_r_169_b : _GEN_12748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12750 = 9'haa == r_count_31_io_out ? io_r_170_b : _GEN_12749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12751 = 9'hab == r_count_31_io_out ? io_r_171_b : _GEN_12750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12752 = 9'hac == r_count_31_io_out ? io_r_172_b : _GEN_12751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12753 = 9'had == r_count_31_io_out ? io_r_173_b : _GEN_12752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12754 = 9'hae == r_count_31_io_out ? io_r_174_b : _GEN_12753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12755 = 9'haf == r_count_31_io_out ? io_r_175_b : _GEN_12754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12756 = 9'hb0 == r_count_31_io_out ? io_r_176_b : _GEN_12755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12757 = 9'hb1 == r_count_31_io_out ? io_r_177_b : _GEN_12756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12758 = 9'hb2 == r_count_31_io_out ? io_r_178_b : _GEN_12757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12759 = 9'hb3 == r_count_31_io_out ? io_r_179_b : _GEN_12758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12760 = 9'hb4 == r_count_31_io_out ? io_r_180_b : _GEN_12759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12761 = 9'hb5 == r_count_31_io_out ? io_r_181_b : _GEN_12760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12762 = 9'hb6 == r_count_31_io_out ? io_r_182_b : _GEN_12761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12763 = 9'hb7 == r_count_31_io_out ? io_r_183_b : _GEN_12762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12764 = 9'hb8 == r_count_31_io_out ? io_r_184_b : _GEN_12763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12765 = 9'hb9 == r_count_31_io_out ? io_r_185_b : _GEN_12764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12766 = 9'hba == r_count_31_io_out ? io_r_186_b : _GEN_12765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12767 = 9'hbb == r_count_31_io_out ? io_r_187_b : _GEN_12766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12768 = 9'hbc == r_count_31_io_out ? io_r_188_b : _GEN_12767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12769 = 9'hbd == r_count_31_io_out ? io_r_189_b : _GEN_12768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12770 = 9'hbe == r_count_31_io_out ? io_r_190_b : _GEN_12769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12771 = 9'hbf == r_count_31_io_out ? io_r_191_b : _GEN_12770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12772 = 9'hc0 == r_count_31_io_out ? io_r_192_b : _GEN_12771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12773 = 9'hc1 == r_count_31_io_out ? io_r_193_b : _GEN_12772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12774 = 9'hc2 == r_count_31_io_out ? io_r_194_b : _GEN_12773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12775 = 9'hc3 == r_count_31_io_out ? io_r_195_b : _GEN_12774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12776 = 9'hc4 == r_count_31_io_out ? io_r_196_b : _GEN_12775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12777 = 9'hc5 == r_count_31_io_out ? io_r_197_b : _GEN_12776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12778 = 9'hc6 == r_count_31_io_out ? io_r_198_b : _GEN_12777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12779 = 9'hc7 == r_count_31_io_out ? io_r_199_b : _GEN_12778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12780 = 9'hc8 == r_count_31_io_out ? io_r_200_b : _GEN_12779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12781 = 9'hc9 == r_count_31_io_out ? io_r_201_b : _GEN_12780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12782 = 9'hca == r_count_31_io_out ? io_r_202_b : _GEN_12781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12783 = 9'hcb == r_count_31_io_out ? io_r_203_b : _GEN_12782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12784 = 9'hcc == r_count_31_io_out ? io_r_204_b : _GEN_12783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12785 = 9'hcd == r_count_31_io_out ? io_r_205_b : _GEN_12784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12786 = 9'hce == r_count_31_io_out ? io_r_206_b : _GEN_12785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12787 = 9'hcf == r_count_31_io_out ? io_r_207_b : _GEN_12786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12788 = 9'hd0 == r_count_31_io_out ? io_r_208_b : _GEN_12787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12789 = 9'hd1 == r_count_31_io_out ? io_r_209_b : _GEN_12788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12790 = 9'hd2 == r_count_31_io_out ? io_r_210_b : _GEN_12789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12791 = 9'hd3 == r_count_31_io_out ? io_r_211_b : _GEN_12790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12792 = 9'hd4 == r_count_31_io_out ? io_r_212_b : _GEN_12791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12793 = 9'hd5 == r_count_31_io_out ? io_r_213_b : _GEN_12792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12794 = 9'hd6 == r_count_31_io_out ? io_r_214_b : _GEN_12793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12795 = 9'hd7 == r_count_31_io_out ? io_r_215_b : _GEN_12794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12796 = 9'hd8 == r_count_31_io_out ? io_r_216_b : _GEN_12795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12797 = 9'hd9 == r_count_31_io_out ? io_r_217_b : _GEN_12796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12798 = 9'hda == r_count_31_io_out ? io_r_218_b : _GEN_12797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12799 = 9'hdb == r_count_31_io_out ? io_r_219_b : _GEN_12798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12800 = 9'hdc == r_count_31_io_out ? io_r_220_b : _GEN_12799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12801 = 9'hdd == r_count_31_io_out ? io_r_221_b : _GEN_12800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12802 = 9'hde == r_count_31_io_out ? io_r_222_b : _GEN_12801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12803 = 9'hdf == r_count_31_io_out ? io_r_223_b : _GEN_12802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12804 = 9'he0 == r_count_31_io_out ? io_r_224_b : _GEN_12803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12805 = 9'he1 == r_count_31_io_out ? io_r_225_b : _GEN_12804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12806 = 9'he2 == r_count_31_io_out ? io_r_226_b : _GEN_12805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12807 = 9'he3 == r_count_31_io_out ? io_r_227_b : _GEN_12806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12808 = 9'he4 == r_count_31_io_out ? io_r_228_b : _GEN_12807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12809 = 9'he5 == r_count_31_io_out ? io_r_229_b : _GEN_12808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12810 = 9'he6 == r_count_31_io_out ? io_r_230_b : _GEN_12809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12811 = 9'he7 == r_count_31_io_out ? io_r_231_b : _GEN_12810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12812 = 9'he8 == r_count_31_io_out ? io_r_232_b : _GEN_12811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12813 = 9'he9 == r_count_31_io_out ? io_r_233_b : _GEN_12812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12814 = 9'hea == r_count_31_io_out ? io_r_234_b : _GEN_12813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12815 = 9'heb == r_count_31_io_out ? io_r_235_b : _GEN_12814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12816 = 9'hec == r_count_31_io_out ? io_r_236_b : _GEN_12815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12817 = 9'hed == r_count_31_io_out ? io_r_237_b : _GEN_12816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12818 = 9'hee == r_count_31_io_out ? io_r_238_b : _GEN_12817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12819 = 9'hef == r_count_31_io_out ? io_r_239_b : _GEN_12818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12820 = 9'hf0 == r_count_31_io_out ? io_r_240_b : _GEN_12819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12821 = 9'hf1 == r_count_31_io_out ? io_r_241_b : _GEN_12820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12822 = 9'hf2 == r_count_31_io_out ? io_r_242_b : _GEN_12821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12823 = 9'hf3 == r_count_31_io_out ? io_r_243_b : _GEN_12822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12824 = 9'hf4 == r_count_31_io_out ? io_r_244_b : _GEN_12823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12825 = 9'hf5 == r_count_31_io_out ? io_r_245_b : _GEN_12824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12826 = 9'hf6 == r_count_31_io_out ? io_r_246_b : _GEN_12825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12827 = 9'hf7 == r_count_31_io_out ? io_r_247_b : _GEN_12826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12828 = 9'hf8 == r_count_31_io_out ? io_r_248_b : _GEN_12827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12829 = 9'hf9 == r_count_31_io_out ? io_r_249_b : _GEN_12828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12830 = 9'hfa == r_count_31_io_out ? io_r_250_b : _GEN_12829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12831 = 9'hfb == r_count_31_io_out ? io_r_251_b : _GEN_12830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12832 = 9'hfc == r_count_31_io_out ? io_r_252_b : _GEN_12831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12833 = 9'hfd == r_count_31_io_out ? io_r_253_b : _GEN_12832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12834 = 9'hfe == r_count_31_io_out ? io_r_254_b : _GEN_12833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12835 = 9'hff == r_count_31_io_out ? io_r_255_b : _GEN_12834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12836 = 9'h100 == r_count_31_io_out ? io_r_256_b : _GEN_12835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12837 = 9'h101 == r_count_31_io_out ? io_r_257_b : _GEN_12836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12838 = 9'h102 == r_count_31_io_out ? io_r_258_b : _GEN_12837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12839 = 9'h103 == r_count_31_io_out ? io_r_259_b : _GEN_12838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12840 = 9'h104 == r_count_31_io_out ? io_r_260_b : _GEN_12839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12841 = 9'h105 == r_count_31_io_out ? io_r_261_b : _GEN_12840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12842 = 9'h106 == r_count_31_io_out ? io_r_262_b : _GEN_12841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12843 = 9'h107 == r_count_31_io_out ? io_r_263_b : _GEN_12842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12844 = 9'h108 == r_count_31_io_out ? io_r_264_b : _GEN_12843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12845 = 9'h109 == r_count_31_io_out ? io_r_265_b : _GEN_12844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12846 = 9'h10a == r_count_31_io_out ? io_r_266_b : _GEN_12845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12847 = 9'h10b == r_count_31_io_out ? io_r_267_b : _GEN_12846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12848 = 9'h10c == r_count_31_io_out ? io_r_268_b : _GEN_12847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12849 = 9'h10d == r_count_31_io_out ? io_r_269_b : _GEN_12848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12850 = 9'h10e == r_count_31_io_out ? io_r_270_b : _GEN_12849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12851 = 9'h10f == r_count_31_io_out ? io_r_271_b : _GEN_12850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12852 = 9'h110 == r_count_31_io_out ? io_r_272_b : _GEN_12851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12853 = 9'h111 == r_count_31_io_out ? io_r_273_b : _GEN_12852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12854 = 9'h112 == r_count_31_io_out ? io_r_274_b : _GEN_12853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12855 = 9'h113 == r_count_31_io_out ? io_r_275_b : _GEN_12854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12856 = 9'h114 == r_count_31_io_out ? io_r_276_b : _GEN_12855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12857 = 9'h115 == r_count_31_io_out ? io_r_277_b : _GEN_12856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12858 = 9'h116 == r_count_31_io_out ? io_r_278_b : _GEN_12857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12859 = 9'h117 == r_count_31_io_out ? io_r_279_b : _GEN_12858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12860 = 9'h118 == r_count_31_io_out ? io_r_280_b : _GEN_12859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12861 = 9'h119 == r_count_31_io_out ? io_r_281_b : _GEN_12860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12862 = 9'h11a == r_count_31_io_out ? io_r_282_b : _GEN_12861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12863 = 9'h11b == r_count_31_io_out ? io_r_283_b : _GEN_12862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12864 = 9'h11c == r_count_31_io_out ? io_r_284_b : _GEN_12863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12865 = 9'h11d == r_count_31_io_out ? io_r_285_b : _GEN_12864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12866 = 9'h11e == r_count_31_io_out ? io_r_286_b : _GEN_12865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12867 = 9'h11f == r_count_31_io_out ? io_r_287_b : _GEN_12866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12868 = 9'h120 == r_count_31_io_out ? io_r_288_b : _GEN_12867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12869 = 9'h121 == r_count_31_io_out ? io_r_289_b : _GEN_12868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12870 = 9'h122 == r_count_31_io_out ? io_r_290_b : _GEN_12869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12871 = 9'h123 == r_count_31_io_out ? io_r_291_b : _GEN_12870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12872 = 9'h124 == r_count_31_io_out ? io_r_292_b : _GEN_12871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12873 = 9'h125 == r_count_31_io_out ? io_r_293_b : _GEN_12872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12874 = 9'h126 == r_count_31_io_out ? io_r_294_b : _GEN_12873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12875 = 9'h127 == r_count_31_io_out ? io_r_295_b : _GEN_12874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12876 = 9'h128 == r_count_31_io_out ? io_r_296_b : _GEN_12875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12877 = 9'h129 == r_count_31_io_out ? io_r_297_b : _GEN_12876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12878 = 9'h12a == r_count_31_io_out ? io_r_298_b : _GEN_12877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12879 = 9'h12b == r_count_31_io_out ? io_r_299_b : _GEN_12878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12880 = 9'h12c == r_count_31_io_out ? io_r_300_b : _GEN_12879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12881 = 9'h12d == r_count_31_io_out ? io_r_301_b : _GEN_12880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12882 = 9'h12e == r_count_31_io_out ? io_r_302_b : _GEN_12881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12883 = 9'h12f == r_count_31_io_out ? io_r_303_b : _GEN_12882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12884 = 9'h130 == r_count_31_io_out ? io_r_304_b : _GEN_12883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12885 = 9'h131 == r_count_31_io_out ? io_r_305_b : _GEN_12884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12886 = 9'h132 == r_count_31_io_out ? io_r_306_b : _GEN_12885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12887 = 9'h133 == r_count_31_io_out ? io_r_307_b : _GEN_12886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12888 = 9'h134 == r_count_31_io_out ? io_r_308_b : _GEN_12887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12889 = 9'h135 == r_count_31_io_out ? io_r_309_b : _GEN_12888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12890 = 9'h136 == r_count_31_io_out ? io_r_310_b : _GEN_12889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12891 = 9'h137 == r_count_31_io_out ? io_r_311_b : _GEN_12890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12892 = 9'h138 == r_count_31_io_out ? io_r_312_b : _GEN_12891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12893 = 9'h139 == r_count_31_io_out ? io_r_313_b : _GEN_12892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12894 = 9'h13a == r_count_31_io_out ? io_r_314_b : _GEN_12893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12895 = 9'h13b == r_count_31_io_out ? io_r_315_b : _GEN_12894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12896 = 9'h13c == r_count_31_io_out ? io_r_316_b : _GEN_12895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12897 = 9'h13d == r_count_31_io_out ? io_r_317_b : _GEN_12896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12898 = 9'h13e == r_count_31_io_out ? io_r_318_b : _GEN_12897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12899 = 9'h13f == r_count_31_io_out ? io_r_319_b : _GEN_12898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12900 = 9'h140 == r_count_31_io_out ? io_r_320_b : _GEN_12899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12901 = 9'h141 == r_count_31_io_out ? io_r_321_b : _GEN_12900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12902 = 9'h142 == r_count_31_io_out ? io_r_322_b : _GEN_12901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12903 = 9'h143 == r_count_31_io_out ? io_r_323_b : _GEN_12902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12904 = 9'h144 == r_count_31_io_out ? io_r_324_b : _GEN_12903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12905 = 9'h145 == r_count_31_io_out ? io_r_325_b : _GEN_12904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12906 = 9'h146 == r_count_31_io_out ? io_r_326_b : _GEN_12905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12907 = 9'h147 == r_count_31_io_out ? io_r_327_b : _GEN_12906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12908 = 9'h148 == r_count_31_io_out ? io_r_328_b : _GEN_12907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12909 = 9'h149 == r_count_31_io_out ? io_r_329_b : _GEN_12908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12910 = 9'h14a == r_count_31_io_out ? io_r_330_b : _GEN_12909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12911 = 9'h14b == r_count_31_io_out ? io_r_331_b : _GEN_12910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12912 = 9'h14c == r_count_31_io_out ? io_r_332_b : _GEN_12911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12913 = 9'h14d == r_count_31_io_out ? io_r_333_b : _GEN_12912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12914 = 9'h14e == r_count_31_io_out ? io_r_334_b : _GEN_12913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12915 = 9'h14f == r_count_31_io_out ? io_r_335_b : _GEN_12914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12916 = 9'h150 == r_count_31_io_out ? io_r_336_b : _GEN_12915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12917 = 9'h151 == r_count_31_io_out ? io_r_337_b : _GEN_12916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12918 = 9'h152 == r_count_31_io_out ? io_r_338_b : _GEN_12917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12919 = 9'h153 == r_count_31_io_out ? io_r_339_b : _GEN_12918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12920 = 9'h154 == r_count_31_io_out ? io_r_340_b : _GEN_12919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12921 = 9'h155 == r_count_31_io_out ? io_r_341_b : _GEN_12920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12922 = 9'h156 == r_count_31_io_out ? io_r_342_b : _GEN_12921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12923 = 9'h157 == r_count_31_io_out ? io_r_343_b : _GEN_12922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12924 = 9'h158 == r_count_31_io_out ? io_r_344_b : _GEN_12923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12925 = 9'h159 == r_count_31_io_out ? io_r_345_b : _GEN_12924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12926 = 9'h15a == r_count_31_io_out ? io_r_346_b : _GEN_12925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12927 = 9'h15b == r_count_31_io_out ? io_r_347_b : _GEN_12926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12928 = 9'h15c == r_count_31_io_out ? io_r_348_b : _GEN_12927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12929 = 9'h15d == r_count_31_io_out ? io_r_349_b : _GEN_12928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12930 = 9'h15e == r_count_31_io_out ? io_r_350_b : _GEN_12929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12931 = 9'h15f == r_count_31_io_out ? io_r_351_b : _GEN_12930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12932 = 9'h160 == r_count_31_io_out ? io_r_352_b : _GEN_12931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12933 = 9'h161 == r_count_31_io_out ? io_r_353_b : _GEN_12932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12934 = 9'h162 == r_count_31_io_out ? io_r_354_b : _GEN_12933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12935 = 9'h163 == r_count_31_io_out ? io_r_355_b : _GEN_12934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12936 = 9'h164 == r_count_31_io_out ? io_r_356_b : _GEN_12935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12937 = 9'h165 == r_count_31_io_out ? io_r_357_b : _GEN_12936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12938 = 9'h166 == r_count_31_io_out ? io_r_358_b : _GEN_12937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12939 = 9'h167 == r_count_31_io_out ? io_r_359_b : _GEN_12938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12940 = 9'h168 == r_count_31_io_out ? io_r_360_b : _GEN_12939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12941 = 9'h169 == r_count_31_io_out ? io_r_361_b : _GEN_12940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12942 = 9'h16a == r_count_31_io_out ? io_r_362_b : _GEN_12941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12943 = 9'h16b == r_count_31_io_out ? io_r_363_b : _GEN_12942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12944 = 9'h16c == r_count_31_io_out ? io_r_364_b : _GEN_12943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12945 = 9'h16d == r_count_31_io_out ? io_r_365_b : _GEN_12944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12946 = 9'h16e == r_count_31_io_out ? io_r_366_b : _GEN_12945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12947 = 9'h16f == r_count_31_io_out ? io_r_367_b : _GEN_12946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12948 = 9'h170 == r_count_31_io_out ? io_r_368_b : _GEN_12947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12949 = 9'h171 == r_count_31_io_out ? io_r_369_b : _GEN_12948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12950 = 9'h172 == r_count_31_io_out ? io_r_370_b : _GEN_12949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12951 = 9'h173 == r_count_31_io_out ? io_r_371_b : _GEN_12950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12952 = 9'h174 == r_count_31_io_out ? io_r_372_b : _GEN_12951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12953 = 9'h175 == r_count_31_io_out ? io_r_373_b : _GEN_12952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12954 = 9'h176 == r_count_31_io_out ? io_r_374_b : _GEN_12953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12955 = 9'h177 == r_count_31_io_out ? io_r_375_b : _GEN_12954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12956 = 9'h178 == r_count_31_io_out ? io_r_376_b : _GEN_12955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12957 = 9'h179 == r_count_31_io_out ? io_r_377_b : _GEN_12956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12958 = 9'h17a == r_count_31_io_out ? io_r_378_b : _GEN_12957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12959 = 9'h17b == r_count_31_io_out ? io_r_379_b : _GEN_12958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12960 = 9'h17c == r_count_31_io_out ? io_r_380_b : _GEN_12959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12961 = 9'h17d == r_count_31_io_out ? io_r_381_b : _GEN_12960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12962 = 9'h17e == r_count_31_io_out ? io_r_382_b : _GEN_12961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12963 = 9'h17f == r_count_31_io_out ? io_r_383_b : _GEN_12962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12964 = 9'h180 == r_count_31_io_out ? io_r_384_b : _GEN_12963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12965 = 9'h181 == r_count_31_io_out ? io_r_385_b : _GEN_12964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12966 = 9'h182 == r_count_31_io_out ? io_r_386_b : _GEN_12965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12967 = 9'h183 == r_count_31_io_out ? io_r_387_b : _GEN_12966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12968 = 9'h184 == r_count_31_io_out ? io_r_388_b : _GEN_12967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12969 = 9'h185 == r_count_31_io_out ? io_r_389_b : _GEN_12968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12970 = 9'h186 == r_count_31_io_out ? io_r_390_b : _GEN_12969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12971 = 9'h187 == r_count_31_io_out ? io_r_391_b : _GEN_12970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12972 = 9'h188 == r_count_31_io_out ? io_r_392_b : _GEN_12971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12973 = 9'h189 == r_count_31_io_out ? io_r_393_b : _GEN_12972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12974 = 9'h18a == r_count_31_io_out ? io_r_394_b : _GEN_12973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12975 = 9'h18b == r_count_31_io_out ? io_r_395_b : _GEN_12974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12976 = 9'h18c == r_count_31_io_out ? io_r_396_b : _GEN_12975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12977 = 9'h18d == r_count_31_io_out ? io_r_397_b : _GEN_12976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12978 = 9'h18e == r_count_31_io_out ? io_r_398_b : _GEN_12977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12981 = 9'h1 == r_count_32_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12982 = 9'h2 == r_count_32_io_out ? io_r_2_b : _GEN_12981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12983 = 9'h3 == r_count_32_io_out ? io_r_3_b : _GEN_12982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12984 = 9'h4 == r_count_32_io_out ? io_r_4_b : _GEN_12983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12985 = 9'h5 == r_count_32_io_out ? io_r_5_b : _GEN_12984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12986 = 9'h6 == r_count_32_io_out ? io_r_6_b : _GEN_12985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12987 = 9'h7 == r_count_32_io_out ? io_r_7_b : _GEN_12986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12988 = 9'h8 == r_count_32_io_out ? io_r_8_b : _GEN_12987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12989 = 9'h9 == r_count_32_io_out ? io_r_9_b : _GEN_12988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12990 = 9'ha == r_count_32_io_out ? io_r_10_b : _GEN_12989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12991 = 9'hb == r_count_32_io_out ? io_r_11_b : _GEN_12990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12992 = 9'hc == r_count_32_io_out ? io_r_12_b : _GEN_12991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12993 = 9'hd == r_count_32_io_out ? io_r_13_b : _GEN_12992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12994 = 9'he == r_count_32_io_out ? io_r_14_b : _GEN_12993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12995 = 9'hf == r_count_32_io_out ? io_r_15_b : _GEN_12994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12996 = 9'h10 == r_count_32_io_out ? io_r_16_b : _GEN_12995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12997 = 9'h11 == r_count_32_io_out ? io_r_17_b : _GEN_12996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12998 = 9'h12 == r_count_32_io_out ? io_r_18_b : _GEN_12997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12999 = 9'h13 == r_count_32_io_out ? io_r_19_b : _GEN_12998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13000 = 9'h14 == r_count_32_io_out ? io_r_20_b : _GEN_12999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13001 = 9'h15 == r_count_32_io_out ? io_r_21_b : _GEN_13000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13002 = 9'h16 == r_count_32_io_out ? io_r_22_b : _GEN_13001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13003 = 9'h17 == r_count_32_io_out ? io_r_23_b : _GEN_13002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13004 = 9'h18 == r_count_32_io_out ? io_r_24_b : _GEN_13003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13005 = 9'h19 == r_count_32_io_out ? io_r_25_b : _GEN_13004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13006 = 9'h1a == r_count_32_io_out ? io_r_26_b : _GEN_13005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13007 = 9'h1b == r_count_32_io_out ? io_r_27_b : _GEN_13006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13008 = 9'h1c == r_count_32_io_out ? io_r_28_b : _GEN_13007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13009 = 9'h1d == r_count_32_io_out ? io_r_29_b : _GEN_13008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13010 = 9'h1e == r_count_32_io_out ? io_r_30_b : _GEN_13009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13011 = 9'h1f == r_count_32_io_out ? io_r_31_b : _GEN_13010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13012 = 9'h20 == r_count_32_io_out ? io_r_32_b : _GEN_13011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13013 = 9'h21 == r_count_32_io_out ? io_r_33_b : _GEN_13012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13014 = 9'h22 == r_count_32_io_out ? io_r_34_b : _GEN_13013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13015 = 9'h23 == r_count_32_io_out ? io_r_35_b : _GEN_13014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13016 = 9'h24 == r_count_32_io_out ? io_r_36_b : _GEN_13015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13017 = 9'h25 == r_count_32_io_out ? io_r_37_b : _GEN_13016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13018 = 9'h26 == r_count_32_io_out ? io_r_38_b : _GEN_13017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13019 = 9'h27 == r_count_32_io_out ? io_r_39_b : _GEN_13018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13020 = 9'h28 == r_count_32_io_out ? io_r_40_b : _GEN_13019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13021 = 9'h29 == r_count_32_io_out ? io_r_41_b : _GEN_13020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13022 = 9'h2a == r_count_32_io_out ? io_r_42_b : _GEN_13021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13023 = 9'h2b == r_count_32_io_out ? io_r_43_b : _GEN_13022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13024 = 9'h2c == r_count_32_io_out ? io_r_44_b : _GEN_13023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13025 = 9'h2d == r_count_32_io_out ? io_r_45_b : _GEN_13024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13026 = 9'h2e == r_count_32_io_out ? io_r_46_b : _GEN_13025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13027 = 9'h2f == r_count_32_io_out ? io_r_47_b : _GEN_13026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13028 = 9'h30 == r_count_32_io_out ? io_r_48_b : _GEN_13027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13029 = 9'h31 == r_count_32_io_out ? io_r_49_b : _GEN_13028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13030 = 9'h32 == r_count_32_io_out ? io_r_50_b : _GEN_13029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13031 = 9'h33 == r_count_32_io_out ? io_r_51_b : _GEN_13030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13032 = 9'h34 == r_count_32_io_out ? io_r_52_b : _GEN_13031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13033 = 9'h35 == r_count_32_io_out ? io_r_53_b : _GEN_13032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13034 = 9'h36 == r_count_32_io_out ? io_r_54_b : _GEN_13033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13035 = 9'h37 == r_count_32_io_out ? io_r_55_b : _GEN_13034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13036 = 9'h38 == r_count_32_io_out ? io_r_56_b : _GEN_13035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13037 = 9'h39 == r_count_32_io_out ? io_r_57_b : _GEN_13036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13038 = 9'h3a == r_count_32_io_out ? io_r_58_b : _GEN_13037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13039 = 9'h3b == r_count_32_io_out ? io_r_59_b : _GEN_13038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13040 = 9'h3c == r_count_32_io_out ? io_r_60_b : _GEN_13039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13041 = 9'h3d == r_count_32_io_out ? io_r_61_b : _GEN_13040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13042 = 9'h3e == r_count_32_io_out ? io_r_62_b : _GEN_13041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13043 = 9'h3f == r_count_32_io_out ? io_r_63_b : _GEN_13042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13044 = 9'h40 == r_count_32_io_out ? io_r_64_b : _GEN_13043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13045 = 9'h41 == r_count_32_io_out ? io_r_65_b : _GEN_13044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13046 = 9'h42 == r_count_32_io_out ? io_r_66_b : _GEN_13045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13047 = 9'h43 == r_count_32_io_out ? io_r_67_b : _GEN_13046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13048 = 9'h44 == r_count_32_io_out ? io_r_68_b : _GEN_13047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13049 = 9'h45 == r_count_32_io_out ? io_r_69_b : _GEN_13048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13050 = 9'h46 == r_count_32_io_out ? io_r_70_b : _GEN_13049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13051 = 9'h47 == r_count_32_io_out ? io_r_71_b : _GEN_13050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13052 = 9'h48 == r_count_32_io_out ? io_r_72_b : _GEN_13051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13053 = 9'h49 == r_count_32_io_out ? io_r_73_b : _GEN_13052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13054 = 9'h4a == r_count_32_io_out ? io_r_74_b : _GEN_13053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13055 = 9'h4b == r_count_32_io_out ? io_r_75_b : _GEN_13054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13056 = 9'h4c == r_count_32_io_out ? io_r_76_b : _GEN_13055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13057 = 9'h4d == r_count_32_io_out ? io_r_77_b : _GEN_13056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13058 = 9'h4e == r_count_32_io_out ? io_r_78_b : _GEN_13057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13059 = 9'h4f == r_count_32_io_out ? io_r_79_b : _GEN_13058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13060 = 9'h50 == r_count_32_io_out ? io_r_80_b : _GEN_13059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13061 = 9'h51 == r_count_32_io_out ? io_r_81_b : _GEN_13060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13062 = 9'h52 == r_count_32_io_out ? io_r_82_b : _GEN_13061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13063 = 9'h53 == r_count_32_io_out ? io_r_83_b : _GEN_13062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13064 = 9'h54 == r_count_32_io_out ? io_r_84_b : _GEN_13063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13065 = 9'h55 == r_count_32_io_out ? io_r_85_b : _GEN_13064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13066 = 9'h56 == r_count_32_io_out ? io_r_86_b : _GEN_13065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13067 = 9'h57 == r_count_32_io_out ? io_r_87_b : _GEN_13066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13068 = 9'h58 == r_count_32_io_out ? io_r_88_b : _GEN_13067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13069 = 9'h59 == r_count_32_io_out ? io_r_89_b : _GEN_13068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13070 = 9'h5a == r_count_32_io_out ? io_r_90_b : _GEN_13069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13071 = 9'h5b == r_count_32_io_out ? io_r_91_b : _GEN_13070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13072 = 9'h5c == r_count_32_io_out ? io_r_92_b : _GEN_13071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13073 = 9'h5d == r_count_32_io_out ? io_r_93_b : _GEN_13072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13074 = 9'h5e == r_count_32_io_out ? io_r_94_b : _GEN_13073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13075 = 9'h5f == r_count_32_io_out ? io_r_95_b : _GEN_13074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13076 = 9'h60 == r_count_32_io_out ? io_r_96_b : _GEN_13075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13077 = 9'h61 == r_count_32_io_out ? io_r_97_b : _GEN_13076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13078 = 9'h62 == r_count_32_io_out ? io_r_98_b : _GEN_13077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13079 = 9'h63 == r_count_32_io_out ? io_r_99_b : _GEN_13078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13080 = 9'h64 == r_count_32_io_out ? io_r_100_b : _GEN_13079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13081 = 9'h65 == r_count_32_io_out ? io_r_101_b : _GEN_13080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13082 = 9'h66 == r_count_32_io_out ? io_r_102_b : _GEN_13081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13083 = 9'h67 == r_count_32_io_out ? io_r_103_b : _GEN_13082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13084 = 9'h68 == r_count_32_io_out ? io_r_104_b : _GEN_13083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13085 = 9'h69 == r_count_32_io_out ? io_r_105_b : _GEN_13084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13086 = 9'h6a == r_count_32_io_out ? io_r_106_b : _GEN_13085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13087 = 9'h6b == r_count_32_io_out ? io_r_107_b : _GEN_13086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13088 = 9'h6c == r_count_32_io_out ? io_r_108_b : _GEN_13087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13089 = 9'h6d == r_count_32_io_out ? io_r_109_b : _GEN_13088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13090 = 9'h6e == r_count_32_io_out ? io_r_110_b : _GEN_13089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13091 = 9'h6f == r_count_32_io_out ? io_r_111_b : _GEN_13090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13092 = 9'h70 == r_count_32_io_out ? io_r_112_b : _GEN_13091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13093 = 9'h71 == r_count_32_io_out ? io_r_113_b : _GEN_13092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13094 = 9'h72 == r_count_32_io_out ? io_r_114_b : _GEN_13093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13095 = 9'h73 == r_count_32_io_out ? io_r_115_b : _GEN_13094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13096 = 9'h74 == r_count_32_io_out ? io_r_116_b : _GEN_13095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13097 = 9'h75 == r_count_32_io_out ? io_r_117_b : _GEN_13096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13098 = 9'h76 == r_count_32_io_out ? io_r_118_b : _GEN_13097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13099 = 9'h77 == r_count_32_io_out ? io_r_119_b : _GEN_13098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13100 = 9'h78 == r_count_32_io_out ? io_r_120_b : _GEN_13099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13101 = 9'h79 == r_count_32_io_out ? io_r_121_b : _GEN_13100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13102 = 9'h7a == r_count_32_io_out ? io_r_122_b : _GEN_13101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13103 = 9'h7b == r_count_32_io_out ? io_r_123_b : _GEN_13102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13104 = 9'h7c == r_count_32_io_out ? io_r_124_b : _GEN_13103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13105 = 9'h7d == r_count_32_io_out ? io_r_125_b : _GEN_13104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13106 = 9'h7e == r_count_32_io_out ? io_r_126_b : _GEN_13105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13107 = 9'h7f == r_count_32_io_out ? io_r_127_b : _GEN_13106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13108 = 9'h80 == r_count_32_io_out ? io_r_128_b : _GEN_13107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13109 = 9'h81 == r_count_32_io_out ? io_r_129_b : _GEN_13108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13110 = 9'h82 == r_count_32_io_out ? io_r_130_b : _GEN_13109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13111 = 9'h83 == r_count_32_io_out ? io_r_131_b : _GEN_13110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13112 = 9'h84 == r_count_32_io_out ? io_r_132_b : _GEN_13111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13113 = 9'h85 == r_count_32_io_out ? io_r_133_b : _GEN_13112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13114 = 9'h86 == r_count_32_io_out ? io_r_134_b : _GEN_13113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13115 = 9'h87 == r_count_32_io_out ? io_r_135_b : _GEN_13114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13116 = 9'h88 == r_count_32_io_out ? io_r_136_b : _GEN_13115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13117 = 9'h89 == r_count_32_io_out ? io_r_137_b : _GEN_13116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13118 = 9'h8a == r_count_32_io_out ? io_r_138_b : _GEN_13117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13119 = 9'h8b == r_count_32_io_out ? io_r_139_b : _GEN_13118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13120 = 9'h8c == r_count_32_io_out ? io_r_140_b : _GEN_13119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13121 = 9'h8d == r_count_32_io_out ? io_r_141_b : _GEN_13120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13122 = 9'h8e == r_count_32_io_out ? io_r_142_b : _GEN_13121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13123 = 9'h8f == r_count_32_io_out ? io_r_143_b : _GEN_13122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13124 = 9'h90 == r_count_32_io_out ? io_r_144_b : _GEN_13123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13125 = 9'h91 == r_count_32_io_out ? io_r_145_b : _GEN_13124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13126 = 9'h92 == r_count_32_io_out ? io_r_146_b : _GEN_13125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13127 = 9'h93 == r_count_32_io_out ? io_r_147_b : _GEN_13126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13128 = 9'h94 == r_count_32_io_out ? io_r_148_b : _GEN_13127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13129 = 9'h95 == r_count_32_io_out ? io_r_149_b : _GEN_13128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13130 = 9'h96 == r_count_32_io_out ? io_r_150_b : _GEN_13129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13131 = 9'h97 == r_count_32_io_out ? io_r_151_b : _GEN_13130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13132 = 9'h98 == r_count_32_io_out ? io_r_152_b : _GEN_13131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13133 = 9'h99 == r_count_32_io_out ? io_r_153_b : _GEN_13132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13134 = 9'h9a == r_count_32_io_out ? io_r_154_b : _GEN_13133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13135 = 9'h9b == r_count_32_io_out ? io_r_155_b : _GEN_13134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13136 = 9'h9c == r_count_32_io_out ? io_r_156_b : _GEN_13135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13137 = 9'h9d == r_count_32_io_out ? io_r_157_b : _GEN_13136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13138 = 9'h9e == r_count_32_io_out ? io_r_158_b : _GEN_13137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13139 = 9'h9f == r_count_32_io_out ? io_r_159_b : _GEN_13138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13140 = 9'ha0 == r_count_32_io_out ? io_r_160_b : _GEN_13139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13141 = 9'ha1 == r_count_32_io_out ? io_r_161_b : _GEN_13140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13142 = 9'ha2 == r_count_32_io_out ? io_r_162_b : _GEN_13141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13143 = 9'ha3 == r_count_32_io_out ? io_r_163_b : _GEN_13142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13144 = 9'ha4 == r_count_32_io_out ? io_r_164_b : _GEN_13143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13145 = 9'ha5 == r_count_32_io_out ? io_r_165_b : _GEN_13144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13146 = 9'ha6 == r_count_32_io_out ? io_r_166_b : _GEN_13145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13147 = 9'ha7 == r_count_32_io_out ? io_r_167_b : _GEN_13146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13148 = 9'ha8 == r_count_32_io_out ? io_r_168_b : _GEN_13147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13149 = 9'ha9 == r_count_32_io_out ? io_r_169_b : _GEN_13148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13150 = 9'haa == r_count_32_io_out ? io_r_170_b : _GEN_13149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13151 = 9'hab == r_count_32_io_out ? io_r_171_b : _GEN_13150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13152 = 9'hac == r_count_32_io_out ? io_r_172_b : _GEN_13151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13153 = 9'had == r_count_32_io_out ? io_r_173_b : _GEN_13152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13154 = 9'hae == r_count_32_io_out ? io_r_174_b : _GEN_13153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13155 = 9'haf == r_count_32_io_out ? io_r_175_b : _GEN_13154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13156 = 9'hb0 == r_count_32_io_out ? io_r_176_b : _GEN_13155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13157 = 9'hb1 == r_count_32_io_out ? io_r_177_b : _GEN_13156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13158 = 9'hb2 == r_count_32_io_out ? io_r_178_b : _GEN_13157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13159 = 9'hb3 == r_count_32_io_out ? io_r_179_b : _GEN_13158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13160 = 9'hb4 == r_count_32_io_out ? io_r_180_b : _GEN_13159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13161 = 9'hb5 == r_count_32_io_out ? io_r_181_b : _GEN_13160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13162 = 9'hb6 == r_count_32_io_out ? io_r_182_b : _GEN_13161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13163 = 9'hb7 == r_count_32_io_out ? io_r_183_b : _GEN_13162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13164 = 9'hb8 == r_count_32_io_out ? io_r_184_b : _GEN_13163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13165 = 9'hb9 == r_count_32_io_out ? io_r_185_b : _GEN_13164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13166 = 9'hba == r_count_32_io_out ? io_r_186_b : _GEN_13165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13167 = 9'hbb == r_count_32_io_out ? io_r_187_b : _GEN_13166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13168 = 9'hbc == r_count_32_io_out ? io_r_188_b : _GEN_13167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13169 = 9'hbd == r_count_32_io_out ? io_r_189_b : _GEN_13168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13170 = 9'hbe == r_count_32_io_out ? io_r_190_b : _GEN_13169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13171 = 9'hbf == r_count_32_io_out ? io_r_191_b : _GEN_13170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13172 = 9'hc0 == r_count_32_io_out ? io_r_192_b : _GEN_13171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13173 = 9'hc1 == r_count_32_io_out ? io_r_193_b : _GEN_13172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13174 = 9'hc2 == r_count_32_io_out ? io_r_194_b : _GEN_13173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13175 = 9'hc3 == r_count_32_io_out ? io_r_195_b : _GEN_13174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13176 = 9'hc4 == r_count_32_io_out ? io_r_196_b : _GEN_13175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13177 = 9'hc5 == r_count_32_io_out ? io_r_197_b : _GEN_13176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13178 = 9'hc6 == r_count_32_io_out ? io_r_198_b : _GEN_13177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13179 = 9'hc7 == r_count_32_io_out ? io_r_199_b : _GEN_13178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13180 = 9'hc8 == r_count_32_io_out ? io_r_200_b : _GEN_13179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13181 = 9'hc9 == r_count_32_io_out ? io_r_201_b : _GEN_13180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13182 = 9'hca == r_count_32_io_out ? io_r_202_b : _GEN_13181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13183 = 9'hcb == r_count_32_io_out ? io_r_203_b : _GEN_13182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13184 = 9'hcc == r_count_32_io_out ? io_r_204_b : _GEN_13183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13185 = 9'hcd == r_count_32_io_out ? io_r_205_b : _GEN_13184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13186 = 9'hce == r_count_32_io_out ? io_r_206_b : _GEN_13185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13187 = 9'hcf == r_count_32_io_out ? io_r_207_b : _GEN_13186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13188 = 9'hd0 == r_count_32_io_out ? io_r_208_b : _GEN_13187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13189 = 9'hd1 == r_count_32_io_out ? io_r_209_b : _GEN_13188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13190 = 9'hd2 == r_count_32_io_out ? io_r_210_b : _GEN_13189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13191 = 9'hd3 == r_count_32_io_out ? io_r_211_b : _GEN_13190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13192 = 9'hd4 == r_count_32_io_out ? io_r_212_b : _GEN_13191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13193 = 9'hd5 == r_count_32_io_out ? io_r_213_b : _GEN_13192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13194 = 9'hd6 == r_count_32_io_out ? io_r_214_b : _GEN_13193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13195 = 9'hd7 == r_count_32_io_out ? io_r_215_b : _GEN_13194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13196 = 9'hd8 == r_count_32_io_out ? io_r_216_b : _GEN_13195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13197 = 9'hd9 == r_count_32_io_out ? io_r_217_b : _GEN_13196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13198 = 9'hda == r_count_32_io_out ? io_r_218_b : _GEN_13197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13199 = 9'hdb == r_count_32_io_out ? io_r_219_b : _GEN_13198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13200 = 9'hdc == r_count_32_io_out ? io_r_220_b : _GEN_13199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13201 = 9'hdd == r_count_32_io_out ? io_r_221_b : _GEN_13200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13202 = 9'hde == r_count_32_io_out ? io_r_222_b : _GEN_13201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13203 = 9'hdf == r_count_32_io_out ? io_r_223_b : _GEN_13202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13204 = 9'he0 == r_count_32_io_out ? io_r_224_b : _GEN_13203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13205 = 9'he1 == r_count_32_io_out ? io_r_225_b : _GEN_13204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13206 = 9'he2 == r_count_32_io_out ? io_r_226_b : _GEN_13205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13207 = 9'he3 == r_count_32_io_out ? io_r_227_b : _GEN_13206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13208 = 9'he4 == r_count_32_io_out ? io_r_228_b : _GEN_13207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13209 = 9'he5 == r_count_32_io_out ? io_r_229_b : _GEN_13208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13210 = 9'he6 == r_count_32_io_out ? io_r_230_b : _GEN_13209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13211 = 9'he7 == r_count_32_io_out ? io_r_231_b : _GEN_13210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13212 = 9'he8 == r_count_32_io_out ? io_r_232_b : _GEN_13211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13213 = 9'he9 == r_count_32_io_out ? io_r_233_b : _GEN_13212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13214 = 9'hea == r_count_32_io_out ? io_r_234_b : _GEN_13213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13215 = 9'heb == r_count_32_io_out ? io_r_235_b : _GEN_13214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13216 = 9'hec == r_count_32_io_out ? io_r_236_b : _GEN_13215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13217 = 9'hed == r_count_32_io_out ? io_r_237_b : _GEN_13216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13218 = 9'hee == r_count_32_io_out ? io_r_238_b : _GEN_13217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13219 = 9'hef == r_count_32_io_out ? io_r_239_b : _GEN_13218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13220 = 9'hf0 == r_count_32_io_out ? io_r_240_b : _GEN_13219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13221 = 9'hf1 == r_count_32_io_out ? io_r_241_b : _GEN_13220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13222 = 9'hf2 == r_count_32_io_out ? io_r_242_b : _GEN_13221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13223 = 9'hf3 == r_count_32_io_out ? io_r_243_b : _GEN_13222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13224 = 9'hf4 == r_count_32_io_out ? io_r_244_b : _GEN_13223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13225 = 9'hf5 == r_count_32_io_out ? io_r_245_b : _GEN_13224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13226 = 9'hf6 == r_count_32_io_out ? io_r_246_b : _GEN_13225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13227 = 9'hf7 == r_count_32_io_out ? io_r_247_b : _GEN_13226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13228 = 9'hf8 == r_count_32_io_out ? io_r_248_b : _GEN_13227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13229 = 9'hf9 == r_count_32_io_out ? io_r_249_b : _GEN_13228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13230 = 9'hfa == r_count_32_io_out ? io_r_250_b : _GEN_13229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13231 = 9'hfb == r_count_32_io_out ? io_r_251_b : _GEN_13230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13232 = 9'hfc == r_count_32_io_out ? io_r_252_b : _GEN_13231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13233 = 9'hfd == r_count_32_io_out ? io_r_253_b : _GEN_13232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13234 = 9'hfe == r_count_32_io_out ? io_r_254_b : _GEN_13233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13235 = 9'hff == r_count_32_io_out ? io_r_255_b : _GEN_13234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13236 = 9'h100 == r_count_32_io_out ? io_r_256_b : _GEN_13235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13237 = 9'h101 == r_count_32_io_out ? io_r_257_b : _GEN_13236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13238 = 9'h102 == r_count_32_io_out ? io_r_258_b : _GEN_13237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13239 = 9'h103 == r_count_32_io_out ? io_r_259_b : _GEN_13238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13240 = 9'h104 == r_count_32_io_out ? io_r_260_b : _GEN_13239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13241 = 9'h105 == r_count_32_io_out ? io_r_261_b : _GEN_13240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13242 = 9'h106 == r_count_32_io_out ? io_r_262_b : _GEN_13241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13243 = 9'h107 == r_count_32_io_out ? io_r_263_b : _GEN_13242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13244 = 9'h108 == r_count_32_io_out ? io_r_264_b : _GEN_13243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13245 = 9'h109 == r_count_32_io_out ? io_r_265_b : _GEN_13244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13246 = 9'h10a == r_count_32_io_out ? io_r_266_b : _GEN_13245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13247 = 9'h10b == r_count_32_io_out ? io_r_267_b : _GEN_13246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13248 = 9'h10c == r_count_32_io_out ? io_r_268_b : _GEN_13247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13249 = 9'h10d == r_count_32_io_out ? io_r_269_b : _GEN_13248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13250 = 9'h10e == r_count_32_io_out ? io_r_270_b : _GEN_13249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13251 = 9'h10f == r_count_32_io_out ? io_r_271_b : _GEN_13250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13252 = 9'h110 == r_count_32_io_out ? io_r_272_b : _GEN_13251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13253 = 9'h111 == r_count_32_io_out ? io_r_273_b : _GEN_13252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13254 = 9'h112 == r_count_32_io_out ? io_r_274_b : _GEN_13253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13255 = 9'h113 == r_count_32_io_out ? io_r_275_b : _GEN_13254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13256 = 9'h114 == r_count_32_io_out ? io_r_276_b : _GEN_13255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13257 = 9'h115 == r_count_32_io_out ? io_r_277_b : _GEN_13256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13258 = 9'h116 == r_count_32_io_out ? io_r_278_b : _GEN_13257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13259 = 9'h117 == r_count_32_io_out ? io_r_279_b : _GEN_13258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13260 = 9'h118 == r_count_32_io_out ? io_r_280_b : _GEN_13259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13261 = 9'h119 == r_count_32_io_out ? io_r_281_b : _GEN_13260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13262 = 9'h11a == r_count_32_io_out ? io_r_282_b : _GEN_13261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13263 = 9'h11b == r_count_32_io_out ? io_r_283_b : _GEN_13262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13264 = 9'h11c == r_count_32_io_out ? io_r_284_b : _GEN_13263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13265 = 9'h11d == r_count_32_io_out ? io_r_285_b : _GEN_13264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13266 = 9'h11e == r_count_32_io_out ? io_r_286_b : _GEN_13265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13267 = 9'h11f == r_count_32_io_out ? io_r_287_b : _GEN_13266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13268 = 9'h120 == r_count_32_io_out ? io_r_288_b : _GEN_13267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13269 = 9'h121 == r_count_32_io_out ? io_r_289_b : _GEN_13268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13270 = 9'h122 == r_count_32_io_out ? io_r_290_b : _GEN_13269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13271 = 9'h123 == r_count_32_io_out ? io_r_291_b : _GEN_13270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13272 = 9'h124 == r_count_32_io_out ? io_r_292_b : _GEN_13271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13273 = 9'h125 == r_count_32_io_out ? io_r_293_b : _GEN_13272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13274 = 9'h126 == r_count_32_io_out ? io_r_294_b : _GEN_13273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13275 = 9'h127 == r_count_32_io_out ? io_r_295_b : _GEN_13274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13276 = 9'h128 == r_count_32_io_out ? io_r_296_b : _GEN_13275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13277 = 9'h129 == r_count_32_io_out ? io_r_297_b : _GEN_13276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13278 = 9'h12a == r_count_32_io_out ? io_r_298_b : _GEN_13277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13279 = 9'h12b == r_count_32_io_out ? io_r_299_b : _GEN_13278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13280 = 9'h12c == r_count_32_io_out ? io_r_300_b : _GEN_13279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13281 = 9'h12d == r_count_32_io_out ? io_r_301_b : _GEN_13280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13282 = 9'h12e == r_count_32_io_out ? io_r_302_b : _GEN_13281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13283 = 9'h12f == r_count_32_io_out ? io_r_303_b : _GEN_13282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13284 = 9'h130 == r_count_32_io_out ? io_r_304_b : _GEN_13283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13285 = 9'h131 == r_count_32_io_out ? io_r_305_b : _GEN_13284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13286 = 9'h132 == r_count_32_io_out ? io_r_306_b : _GEN_13285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13287 = 9'h133 == r_count_32_io_out ? io_r_307_b : _GEN_13286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13288 = 9'h134 == r_count_32_io_out ? io_r_308_b : _GEN_13287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13289 = 9'h135 == r_count_32_io_out ? io_r_309_b : _GEN_13288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13290 = 9'h136 == r_count_32_io_out ? io_r_310_b : _GEN_13289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13291 = 9'h137 == r_count_32_io_out ? io_r_311_b : _GEN_13290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13292 = 9'h138 == r_count_32_io_out ? io_r_312_b : _GEN_13291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13293 = 9'h139 == r_count_32_io_out ? io_r_313_b : _GEN_13292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13294 = 9'h13a == r_count_32_io_out ? io_r_314_b : _GEN_13293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13295 = 9'h13b == r_count_32_io_out ? io_r_315_b : _GEN_13294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13296 = 9'h13c == r_count_32_io_out ? io_r_316_b : _GEN_13295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13297 = 9'h13d == r_count_32_io_out ? io_r_317_b : _GEN_13296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13298 = 9'h13e == r_count_32_io_out ? io_r_318_b : _GEN_13297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13299 = 9'h13f == r_count_32_io_out ? io_r_319_b : _GEN_13298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13300 = 9'h140 == r_count_32_io_out ? io_r_320_b : _GEN_13299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13301 = 9'h141 == r_count_32_io_out ? io_r_321_b : _GEN_13300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13302 = 9'h142 == r_count_32_io_out ? io_r_322_b : _GEN_13301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13303 = 9'h143 == r_count_32_io_out ? io_r_323_b : _GEN_13302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13304 = 9'h144 == r_count_32_io_out ? io_r_324_b : _GEN_13303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13305 = 9'h145 == r_count_32_io_out ? io_r_325_b : _GEN_13304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13306 = 9'h146 == r_count_32_io_out ? io_r_326_b : _GEN_13305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13307 = 9'h147 == r_count_32_io_out ? io_r_327_b : _GEN_13306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13308 = 9'h148 == r_count_32_io_out ? io_r_328_b : _GEN_13307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13309 = 9'h149 == r_count_32_io_out ? io_r_329_b : _GEN_13308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13310 = 9'h14a == r_count_32_io_out ? io_r_330_b : _GEN_13309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13311 = 9'h14b == r_count_32_io_out ? io_r_331_b : _GEN_13310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13312 = 9'h14c == r_count_32_io_out ? io_r_332_b : _GEN_13311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13313 = 9'h14d == r_count_32_io_out ? io_r_333_b : _GEN_13312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13314 = 9'h14e == r_count_32_io_out ? io_r_334_b : _GEN_13313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13315 = 9'h14f == r_count_32_io_out ? io_r_335_b : _GEN_13314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13316 = 9'h150 == r_count_32_io_out ? io_r_336_b : _GEN_13315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13317 = 9'h151 == r_count_32_io_out ? io_r_337_b : _GEN_13316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13318 = 9'h152 == r_count_32_io_out ? io_r_338_b : _GEN_13317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13319 = 9'h153 == r_count_32_io_out ? io_r_339_b : _GEN_13318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13320 = 9'h154 == r_count_32_io_out ? io_r_340_b : _GEN_13319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13321 = 9'h155 == r_count_32_io_out ? io_r_341_b : _GEN_13320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13322 = 9'h156 == r_count_32_io_out ? io_r_342_b : _GEN_13321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13323 = 9'h157 == r_count_32_io_out ? io_r_343_b : _GEN_13322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13324 = 9'h158 == r_count_32_io_out ? io_r_344_b : _GEN_13323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13325 = 9'h159 == r_count_32_io_out ? io_r_345_b : _GEN_13324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13326 = 9'h15a == r_count_32_io_out ? io_r_346_b : _GEN_13325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13327 = 9'h15b == r_count_32_io_out ? io_r_347_b : _GEN_13326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13328 = 9'h15c == r_count_32_io_out ? io_r_348_b : _GEN_13327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13329 = 9'h15d == r_count_32_io_out ? io_r_349_b : _GEN_13328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13330 = 9'h15e == r_count_32_io_out ? io_r_350_b : _GEN_13329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13331 = 9'h15f == r_count_32_io_out ? io_r_351_b : _GEN_13330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13332 = 9'h160 == r_count_32_io_out ? io_r_352_b : _GEN_13331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13333 = 9'h161 == r_count_32_io_out ? io_r_353_b : _GEN_13332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13334 = 9'h162 == r_count_32_io_out ? io_r_354_b : _GEN_13333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13335 = 9'h163 == r_count_32_io_out ? io_r_355_b : _GEN_13334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13336 = 9'h164 == r_count_32_io_out ? io_r_356_b : _GEN_13335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13337 = 9'h165 == r_count_32_io_out ? io_r_357_b : _GEN_13336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13338 = 9'h166 == r_count_32_io_out ? io_r_358_b : _GEN_13337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13339 = 9'h167 == r_count_32_io_out ? io_r_359_b : _GEN_13338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13340 = 9'h168 == r_count_32_io_out ? io_r_360_b : _GEN_13339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13341 = 9'h169 == r_count_32_io_out ? io_r_361_b : _GEN_13340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13342 = 9'h16a == r_count_32_io_out ? io_r_362_b : _GEN_13341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13343 = 9'h16b == r_count_32_io_out ? io_r_363_b : _GEN_13342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13344 = 9'h16c == r_count_32_io_out ? io_r_364_b : _GEN_13343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13345 = 9'h16d == r_count_32_io_out ? io_r_365_b : _GEN_13344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13346 = 9'h16e == r_count_32_io_out ? io_r_366_b : _GEN_13345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13347 = 9'h16f == r_count_32_io_out ? io_r_367_b : _GEN_13346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13348 = 9'h170 == r_count_32_io_out ? io_r_368_b : _GEN_13347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13349 = 9'h171 == r_count_32_io_out ? io_r_369_b : _GEN_13348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13350 = 9'h172 == r_count_32_io_out ? io_r_370_b : _GEN_13349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13351 = 9'h173 == r_count_32_io_out ? io_r_371_b : _GEN_13350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13352 = 9'h174 == r_count_32_io_out ? io_r_372_b : _GEN_13351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13353 = 9'h175 == r_count_32_io_out ? io_r_373_b : _GEN_13352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13354 = 9'h176 == r_count_32_io_out ? io_r_374_b : _GEN_13353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13355 = 9'h177 == r_count_32_io_out ? io_r_375_b : _GEN_13354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13356 = 9'h178 == r_count_32_io_out ? io_r_376_b : _GEN_13355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13357 = 9'h179 == r_count_32_io_out ? io_r_377_b : _GEN_13356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13358 = 9'h17a == r_count_32_io_out ? io_r_378_b : _GEN_13357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13359 = 9'h17b == r_count_32_io_out ? io_r_379_b : _GEN_13358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13360 = 9'h17c == r_count_32_io_out ? io_r_380_b : _GEN_13359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13361 = 9'h17d == r_count_32_io_out ? io_r_381_b : _GEN_13360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13362 = 9'h17e == r_count_32_io_out ? io_r_382_b : _GEN_13361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13363 = 9'h17f == r_count_32_io_out ? io_r_383_b : _GEN_13362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13364 = 9'h180 == r_count_32_io_out ? io_r_384_b : _GEN_13363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13365 = 9'h181 == r_count_32_io_out ? io_r_385_b : _GEN_13364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13366 = 9'h182 == r_count_32_io_out ? io_r_386_b : _GEN_13365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13367 = 9'h183 == r_count_32_io_out ? io_r_387_b : _GEN_13366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13368 = 9'h184 == r_count_32_io_out ? io_r_388_b : _GEN_13367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13369 = 9'h185 == r_count_32_io_out ? io_r_389_b : _GEN_13368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13370 = 9'h186 == r_count_32_io_out ? io_r_390_b : _GEN_13369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13371 = 9'h187 == r_count_32_io_out ? io_r_391_b : _GEN_13370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13372 = 9'h188 == r_count_32_io_out ? io_r_392_b : _GEN_13371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13373 = 9'h189 == r_count_32_io_out ? io_r_393_b : _GEN_13372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13374 = 9'h18a == r_count_32_io_out ? io_r_394_b : _GEN_13373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13375 = 9'h18b == r_count_32_io_out ? io_r_395_b : _GEN_13374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13376 = 9'h18c == r_count_32_io_out ? io_r_396_b : _GEN_13375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13377 = 9'h18d == r_count_32_io_out ? io_r_397_b : _GEN_13376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13378 = 9'h18e == r_count_32_io_out ? io_r_398_b : _GEN_13377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13381 = 9'h1 == r_count_33_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13382 = 9'h2 == r_count_33_io_out ? io_r_2_b : _GEN_13381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13383 = 9'h3 == r_count_33_io_out ? io_r_3_b : _GEN_13382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13384 = 9'h4 == r_count_33_io_out ? io_r_4_b : _GEN_13383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13385 = 9'h5 == r_count_33_io_out ? io_r_5_b : _GEN_13384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13386 = 9'h6 == r_count_33_io_out ? io_r_6_b : _GEN_13385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13387 = 9'h7 == r_count_33_io_out ? io_r_7_b : _GEN_13386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13388 = 9'h8 == r_count_33_io_out ? io_r_8_b : _GEN_13387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13389 = 9'h9 == r_count_33_io_out ? io_r_9_b : _GEN_13388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13390 = 9'ha == r_count_33_io_out ? io_r_10_b : _GEN_13389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13391 = 9'hb == r_count_33_io_out ? io_r_11_b : _GEN_13390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13392 = 9'hc == r_count_33_io_out ? io_r_12_b : _GEN_13391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13393 = 9'hd == r_count_33_io_out ? io_r_13_b : _GEN_13392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13394 = 9'he == r_count_33_io_out ? io_r_14_b : _GEN_13393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13395 = 9'hf == r_count_33_io_out ? io_r_15_b : _GEN_13394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13396 = 9'h10 == r_count_33_io_out ? io_r_16_b : _GEN_13395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13397 = 9'h11 == r_count_33_io_out ? io_r_17_b : _GEN_13396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13398 = 9'h12 == r_count_33_io_out ? io_r_18_b : _GEN_13397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13399 = 9'h13 == r_count_33_io_out ? io_r_19_b : _GEN_13398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13400 = 9'h14 == r_count_33_io_out ? io_r_20_b : _GEN_13399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13401 = 9'h15 == r_count_33_io_out ? io_r_21_b : _GEN_13400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13402 = 9'h16 == r_count_33_io_out ? io_r_22_b : _GEN_13401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13403 = 9'h17 == r_count_33_io_out ? io_r_23_b : _GEN_13402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13404 = 9'h18 == r_count_33_io_out ? io_r_24_b : _GEN_13403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13405 = 9'h19 == r_count_33_io_out ? io_r_25_b : _GEN_13404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13406 = 9'h1a == r_count_33_io_out ? io_r_26_b : _GEN_13405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13407 = 9'h1b == r_count_33_io_out ? io_r_27_b : _GEN_13406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13408 = 9'h1c == r_count_33_io_out ? io_r_28_b : _GEN_13407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13409 = 9'h1d == r_count_33_io_out ? io_r_29_b : _GEN_13408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13410 = 9'h1e == r_count_33_io_out ? io_r_30_b : _GEN_13409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13411 = 9'h1f == r_count_33_io_out ? io_r_31_b : _GEN_13410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13412 = 9'h20 == r_count_33_io_out ? io_r_32_b : _GEN_13411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13413 = 9'h21 == r_count_33_io_out ? io_r_33_b : _GEN_13412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13414 = 9'h22 == r_count_33_io_out ? io_r_34_b : _GEN_13413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13415 = 9'h23 == r_count_33_io_out ? io_r_35_b : _GEN_13414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13416 = 9'h24 == r_count_33_io_out ? io_r_36_b : _GEN_13415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13417 = 9'h25 == r_count_33_io_out ? io_r_37_b : _GEN_13416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13418 = 9'h26 == r_count_33_io_out ? io_r_38_b : _GEN_13417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13419 = 9'h27 == r_count_33_io_out ? io_r_39_b : _GEN_13418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13420 = 9'h28 == r_count_33_io_out ? io_r_40_b : _GEN_13419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13421 = 9'h29 == r_count_33_io_out ? io_r_41_b : _GEN_13420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13422 = 9'h2a == r_count_33_io_out ? io_r_42_b : _GEN_13421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13423 = 9'h2b == r_count_33_io_out ? io_r_43_b : _GEN_13422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13424 = 9'h2c == r_count_33_io_out ? io_r_44_b : _GEN_13423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13425 = 9'h2d == r_count_33_io_out ? io_r_45_b : _GEN_13424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13426 = 9'h2e == r_count_33_io_out ? io_r_46_b : _GEN_13425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13427 = 9'h2f == r_count_33_io_out ? io_r_47_b : _GEN_13426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13428 = 9'h30 == r_count_33_io_out ? io_r_48_b : _GEN_13427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13429 = 9'h31 == r_count_33_io_out ? io_r_49_b : _GEN_13428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13430 = 9'h32 == r_count_33_io_out ? io_r_50_b : _GEN_13429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13431 = 9'h33 == r_count_33_io_out ? io_r_51_b : _GEN_13430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13432 = 9'h34 == r_count_33_io_out ? io_r_52_b : _GEN_13431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13433 = 9'h35 == r_count_33_io_out ? io_r_53_b : _GEN_13432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13434 = 9'h36 == r_count_33_io_out ? io_r_54_b : _GEN_13433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13435 = 9'h37 == r_count_33_io_out ? io_r_55_b : _GEN_13434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13436 = 9'h38 == r_count_33_io_out ? io_r_56_b : _GEN_13435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13437 = 9'h39 == r_count_33_io_out ? io_r_57_b : _GEN_13436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13438 = 9'h3a == r_count_33_io_out ? io_r_58_b : _GEN_13437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13439 = 9'h3b == r_count_33_io_out ? io_r_59_b : _GEN_13438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13440 = 9'h3c == r_count_33_io_out ? io_r_60_b : _GEN_13439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13441 = 9'h3d == r_count_33_io_out ? io_r_61_b : _GEN_13440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13442 = 9'h3e == r_count_33_io_out ? io_r_62_b : _GEN_13441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13443 = 9'h3f == r_count_33_io_out ? io_r_63_b : _GEN_13442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13444 = 9'h40 == r_count_33_io_out ? io_r_64_b : _GEN_13443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13445 = 9'h41 == r_count_33_io_out ? io_r_65_b : _GEN_13444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13446 = 9'h42 == r_count_33_io_out ? io_r_66_b : _GEN_13445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13447 = 9'h43 == r_count_33_io_out ? io_r_67_b : _GEN_13446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13448 = 9'h44 == r_count_33_io_out ? io_r_68_b : _GEN_13447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13449 = 9'h45 == r_count_33_io_out ? io_r_69_b : _GEN_13448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13450 = 9'h46 == r_count_33_io_out ? io_r_70_b : _GEN_13449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13451 = 9'h47 == r_count_33_io_out ? io_r_71_b : _GEN_13450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13452 = 9'h48 == r_count_33_io_out ? io_r_72_b : _GEN_13451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13453 = 9'h49 == r_count_33_io_out ? io_r_73_b : _GEN_13452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13454 = 9'h4a == r_count_33_io_out ? io_r_74_b : _GEN_13453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13455 = 9'h4b == r_count_33_io_out ? io_r_75_b : _GEN_13454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13456 = 9'h4c == r_count_33_io_out ? io_r_76_b : _GEN_13455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13457 = 9'h4d == r_count_33_io_out ? io_r_77_b : _GEN_13456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13458 = 9'h4e == r_count_33_io_out ? io_r_78_b : _GEN_13457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13459 = 9'h4f == r_count_33_io_out ? io_r_79_b : _GEN_13458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13460 = 9'h50 == r_count_33_io_out ? io_r_80_b : _GEN_13459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13461 = 9'h51 == r_count_33_io_out ? io_r_81_b : _GEN_13460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13462 = 9'h52 == r_count_33_io_out ? io_r_82_b : _GEN_13461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13463 = 9'h53 == r_count_33_io_out ? io_r_83_b : _GEN_13462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13464 = 9'h54 == r_count_33_io_out ? io_r_84_b : _GEN_13463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13465 = 9'h55 == r_count_33_io_out ? io_r_85_b : _GEN_13464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13466 = 9'h56 == r_count_33_io_out ? io_r_86_b : _GEN_13465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13467 = 9'h57 == r_count_33_io_out ? io_r_87_b : _GEN_13466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13468 = 9'h58 == r_count_33_io_out ? io_r_88_b : _GEN_13467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13469 = 9'h59 == r_count_33_io_out ? io_r_89_b : _GEN_13468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13470 = 9'h5a == r_count_33_io_out ? io_r_90_b : _GEN_13469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13471 = 9'h5b == r_count_33_io_out ? io_r_91_b : _GEN_13470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13472 = 9'h5c == r_count_33_io_out ? io_r_92_b : _GEN_13471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13473 = 9'h5d == r_count_33_io_out ? io_r_93_b : _GEN_13472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13474 = 9'h5e == r_count_33_io_out ? io_r_94_b : _GEN_13473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13475 = 9'h5f == r_count_33_io_out ? io_r_95_b : _GEN_13474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13476 = 9'h60 == r_count_33_io_out ? io_r_96_b : _GEN_13475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13477 = 9'h61 == r_count_33_io_out ? io_r_97_b : _GEN_13476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13478 = 9'h62 == r_count_33_io_out ? io_r_98_b : _GEN_13477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13479 = 9'h63 == r_count_33_io_out ? io_r_99_b : _GEN_13478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13480 = 9'h64 == r_count_33_io_out ? io_r_100_b : _GEN_13479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13481 = 9'h65 == r_count_33_io_out ? io_r_101_b : _GEN_13480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13482 = 9'h66 == r_count_33_io_out ? io_r_102_b : _GEN_13481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13483 = 9'h67 == r_count_33_io_out ? io_r_103_b : _GEN_13482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13484 = 9'h68 == r_count_33_io_out ? io_r_104_b : _GEN_13483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13485 = 9'h69 == r_count_33_io_out ? io_r_105_b : _GEN_13484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13486 = 9'h6a == r_count_33_io_out ? io_r_106_b : _GEN_13485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13487 = 9'h6b == r_count_33_io_out ? io_r_107_b : _GEN_13486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13488 = 9'h6c == r_count_33_io_out ? io_r_108_b : _GEN_13487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13489 = 9'h6d == r_count_33_io_out ? io_r_109_b : _GEN_13488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13490 = 9'h6e == r_count_33_io_out ? io_r_110_b : _GEN_13489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13491 = 9'h6f == r_count_33_io_out ? io_r_111_b : _GEN_13490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13492 = 9'h70 == r_count_33_io_out ? io_r_112_b : _GEN_13491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13493 = 9'h71 == r_count_33_io_out ? io_r_113_b : _GEN_13492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13494 = 9'h72 == r_count_33_io_out ? io_r_114_b : _GEN_13493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13495 = 9'h73 == r_count_33_io_out ? io_r_115_b : _GEN_13494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13496 = 9'h74 == r_count_33_io_out ? io_r_116_b : _GEN_13495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13497 = 9'h75 == r_count_33_io_out ? io_r_117_b : _GEN_13496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13498 = 9'h76 == r_count_33_io_out ? io_r_118_b : _GEN_13497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13499 = 9'h77 == r_count_33_io_out ? io_r_119_b : _GEN_13498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13500 = 9'h78 == r_count_33_io_out ? io_r_120_b : _GEN_13499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13501 = 9'h79 == r_count_33_io_out ? io_r_121_b : _GEN_13500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13502 = 9'h7a == r_count_33_io_out ? io_r_122_b : _GEN_13501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13503 = 9'h7b == r_count_33_io_out ? io_r_123_b : _GEN_13502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13504 = 9'h7c == r_count_33_io_out ? io_r_124_b : _GEN_13503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13505 = 9'h7d == r_count_33_io_out ? io_r_125_b : _GEN_13504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13506 = 9'h7e == r_count_33_io_out ? io_r_126_b : _GEN_13505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13507 = 9'h7f == r_count_33_io_out ? io_r_127_b : _GEN_13506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13508 = 9'h80 == r_count_33_io_out ? io_r_128_b : _GEN_13507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13509 = 9'h81 == r_count_33_io_out ? io_r_129_b : _GEN_13508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13510 = 9'h82 == r_count_33_io_out ? io_r_130_b : _GEN_13509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13511 = 9'h83 == r_count_33_io_out ? io_r_131_b : _GEN_13510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13512 = 9'h84 == r_count_33_io_out ? io_r_132_b : _GEN_13511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13513 = 9'h85 == r_count_33_io_out ? io_r_133_b : _GEN_13512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13514 = 9'h86 == r_count_33_io_out ? io_r_134_b : _GEN_13513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13515 = 9'h87 == r_count_33_io_out ? io_r_135_b : _GEN_13514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13516 = 9'h88 == r_count_33_io_out ? io_r_136_b : _GEN_13515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13517 = 9'h89 == r_count_33_io_out ? io_r_137_b : _GEN_13516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13518 = 9'h8a == r_count_33_io_out ? io_r_138_b : _GEN_13517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13519 = 9'h8b == r_count_33_io_out ? io_r_139_b : _GEN_13518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13520 = 9'h8c == r_count_33_io_out ? io_r_140_b : _GEN_13519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13521 = 9'h8d == r_count_33_io_out ? io_r_141_b : _GEN_13520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13522 = 9'h8e == r_count_33_io_out ? io_r_142_b : _GEN_13521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13523 = 9'h8f == r_count_33_io_out ? io_r_143_b : _GEN_13522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13524 = 9'h90 == r_count_33_io_out ? io_r_144_b : _GEN_13523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13525 = 9'h91 == r_count_33_io_out ? io_r_145_b : _GEN_13524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13526 = 9'h92 == r_count_33_io_out ? io_r_146_b : _GEN_13525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13527 = 9'h93 == r_count_33_io_out ? io_r_147_b : _GEN_13526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13528 = 9'h94 == r_count_33_io_out ? io_r_148_b : _GEN_13527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13529 = 9'h95 == r_count_33_io_out ? io_r_149_b : _GEN_13528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13530 = 9'h96 == r_count_33_io_out ? io_r_150_b : _GEN_13529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13531 = 9'h97 == r_count_33_io_out ? io_r_151_b : _GEN_13530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13532 = 9'h98 == r_count_33_io_out ? io_r_152_b : _GEN_13531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13533 = 9'h99 == r_count_33_io_out ? io_r_153_b : _GEN_13532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13534 = 9'h9a == r_count_33_io_out ? io_r_154_b : _GEN_13533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13535 = 9'h9b == r_count_33_io_out ? io_r_155_b : _GEN_13534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13536 = 9'h9c == r_count_33_io_out ? io_r_156_b : _GEN_13535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13537 = 9'h9d == r_count_33_io_out ? io_r_157_b : _GEN_13536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13538 = 9'h9e == r_count_33_io_out ? io_r_158_b : _GEN_13537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13539 = 9'h9f == r_count_33_io_out ? io_r_159_b : _GEN_13538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13540 = 9'ha0 == r_count_33_io_out ? io_r_160_b : _GEN_13539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13541 = 9'ha1 == r_count_33_io_out ? io_r_161_b : _GEN_13540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13542 = 9'ha2 == r_count_33_io_out ? io_r_162_b : _GEN_13541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13543 = 9'ha3 == r_count_33_io_out ? io_r_163_b : _GEN_13542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13544 = 9'ha4 == r_count_33_io_out ? io_r_164_b : _GEN_13543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13545 = 9'ha5 == r_count_33_io_out ? io_r_165_b : _GEN_13544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13546 = 9'ha6 == r_count_33_io_out ? io_r_166_b : _GEN_13545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13547 = 9'ha7 == r_count_33_io_out ? io_r_167_b : _GEN_13546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13548 = 9'ha8 == r_count_33_io_out ? io_r_168_b : _GEN_13547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13549 = 9'ha9 == r_count_33_io_out ? io_r_169_b : _GEN_13548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13550 = 9'haa == r_count_33_io_out ? io_r_170_b : _GEN_13549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13551 = 9'hab == r_count_33_io_out ? io_r_171_b : _GEN_13550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13552 = 9'hac == r_count_33_io_out ? io_r_172_b : _GEN_13551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13553 = 9'had == r_count_33_io_out ? io_r_173_b : _GEN_13552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13554 = 9'hae == r_count_33_io_out ? io_r_174_b : _GEN_13553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13555 = 9'haf == r_count_33_io_out ? io_r_175_b : _GEN_13554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13556 = 9'hb0 == r_count_33_io_out ? io_r_176_b : _GEN_13555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13557 = 9'hb1 == r_count_33_io_out ? io_r_177_b : _GEN_13556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13558 = 9'hb2 == r_count_33_io_out ? io_r_178_b : _GEN_13557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13559 = 9'hb3 == r_count_33_io_out ? io_r_179_b : _GEN_13558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13560 = 9'hb4 == r_count_33_io_out ? io_r_180_b : _GEN_13559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13561 = 9'hb5 == r_count_33_io_out ? io_r_181_b : _GEN_13560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13562 = 9'hb6 == r_count_33_io_out ? io_r_182_b : _GEN_13561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13563 = 9'hb7 == r_count_33_io_out ? io_r_183_b : _GEN_13562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13564 = 9'hb8 == r_count_33_io_out ? io_r_184_b : _GEN_13563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13565 = 9'hb9 == r_count_33_io_out ? io_r_185_b : _GEN_13564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13566 = 9'hba == r_count_33_io_out ? io_r_186_b : _GEN_13565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13567 = 9'hbb == r_count_33_io_out ? io_r_187_b : _GEN_13566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13568 = 9'hbc == r_count_33_io_out ? io_r_188_b : _GEN_13567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13569 = 9'hbd == r_count_33_io_out ? io_r_189_b : _GEN_13568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13570 = 9'hbe == r_count_33_io_out ? io_r_190_b : _GEN_13569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13571 = 9'hbf == r_count_33_io_out ? io_r_191_b : _GEN_13570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13572 = 9'hc0 == r_count_33_io_out ? io_r_192_b : _GEN_13571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13573 = 9'hc1 == r_count_33_io_out ? io_r_193_b : _GEN_13572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13574 = 9'hc2 == r_count_33_io_out ? io_r_194_b : _GEN_13573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13575 = 9'hc3 == r_count_33_io_out ? io_r_195_b : _GEN_13574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13576 = 9'hc4 == r_count_33_io_out ? io_r_196_b : _GEN_13575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13577 = 9'hc5 == r_count_33_io_out ? io_r_197_b : _GEN_13576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13578 = 9'hc6 == r_count_33_io_out ? io_r_198_b : _GEN_13577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13579 = 9'hc7 == r_count_33_io_out ? io_r_199_b : _GEN_13578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13580 = 9'hc8 == r_count_33_io_out ? io_r_200_b : _GEN_13579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13581 = 9'hc9 == r_count_33_io_out ? io_r_201_b : _GEN_13580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13582 = 9'hca == r_count_33_io_out ? io_r_202_b : _GEN_13581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13583 = 9'hcb == r_count_33_io_out ? io_r_203_b : _GEN_13582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13584 = 9'hcc == r_count_33_io_out ? io_r_204_b : _GEN_13583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13585 = 9'hcd == r_count_33_io_out ? io_r_205_b : _GEN_13584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13586 = 9'hce == r_count_33_io_out ? io_r_206_b : _GEN_13585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13587 = 9'hcf == r_count_33_io_out ? io_r_207_b : _GEN_13586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13588 = 9'hd0 == r_count_33_io_out ? io_r_208_b : _GEN_13587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13589 = 9'hd1 == r_count_33_io_out ? io_r_209_b : _GEN_13588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13590 = 9'hd2 == r_count_33_io_out ? io_r_210_b : _GEN_13589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13591 = 9'hd3 == r_count_33_io_out ? io_r_211_b : _GEN_13590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13592 = 9'hd4 == r_count_33_io_out ? io_r_212_b : _GEN_13591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13593 = 9'hd5 == r_count_33_io_out ? io_r_213_b : _GEN_13592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13594 = 9'hd6 == r_count_33_io_out ? io_r_214_b : _GEN_13593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13595 = 9'hd7 == r_count_33_io_out ? io_r_215_b : _GEN_13594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13596 = 9'hd8 == r_count_33_io_out ? io_r_216_b : _GEN_13595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13597 = 9'hd9 == r_count_33_io_out ? io_r_217_b : _GEN_13596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13598 = 9'hda == r_count_33_io_out ? io_r_218_b : _GEN_13597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13599 = 9'hdb == r_count_33_io_out ? io_r_219_b : _GEN_13598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13600 = 9'hdc == r_count_33_io_out ? io_r_220_b : _GEN_13599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13601 = 9'hdd == r_count_33_io_out ? io_r_221_b : _GEN_13600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13602 = 9'hde == r_count_33_io_out ? io_r_222_b : _GEN_13601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13603 = 9'hdf == r_count_33_io_out ? io_r_223_b : _GEN_13602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13604 = 9'he0 == r_count_33_io_out ? io_r_224_b : _GEN_13603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13605 = 9'he1 == r_count_33_io_out ? io_r_225_b : _GEN_13604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13606 = 9'he2 == r_count_33_io_out ? io_r_226_b : _GEN_13605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13607 = 9'he3 == r_count_33_io_out ? io_r_227_b : _GEN_13606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13608 = 9'he4 == r_count_33_io_out ? io_r_228_b : _GEN_13607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13609 = 9'he5 == r_count_33_io_out ? io_r_229_b : _GEN_13608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13610 = 9'he6 == r_count_33_io_out ? io_r_230_b : _GEN_13609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13611 = 9'he7 == r_count_33_io_out ? io_r_231_b : _GEN_13610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13612 = 9'he8 == r_count_33_io_out ? io_r_232_b : _GEN_13611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13613 = 9'he9 == r_count_33_io_out ? io_r_233_b : _GEN_13612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13614 = 9'hea == r_count_33_io_out ? io_r_234_b : _GEN_13613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13615 = 9'heb == r_count_33_io_out ? io_r_235_b : _GEN_13614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13616 = 9'hec == r_count_33_io_out ? io_r_236_b : _GEN_13615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13617 = 9'hed == r_count_33_io_out ? io_r_237_b : _GEN_13616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13618 = 9'hee == r_count_33_io_out ? io_r_238_b : _GEN_13617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13619 = 9'hef == r_count_33_io_out ? io_r_239_b : _GEN_13618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13620 = 9'hf0 == r_count_33_io_out ? io_r_240_b : _GEN_13619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13621 = 9'hf1 == r_count_33_io_out ? io_r_241_b : _GEN_13620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13622 = 9'hf2 == r_count_33_io_out ? io_r_242_b : _GEN_13621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13623 = 9'hf3 == r_count_33_io_out ? io_r_243_b : _GEN_13622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13624 = 9'hf4 == r_count_33_io_out ? io_r_244_b : _GEN_13623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13625 = 9'hf5 == r_count_33_io_out ? io_r_245_b : _GEN_13624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13626 = 9'hf6 == r_count_33_io_out ? io_r_246_b : _GEN_13625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13627 = 9'hf7 == r_count_33_io_out ? io_r_247_b : _GEN_13626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13628 = 9'hf8 == r_count_33_io_out ? io_r_248_b : _GEN_13627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13629 = 9'hf9 == r_count_33_io_out ? io_r_249_b : _GEN_13628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13630 = 9'hfa == r_count_33_io_out ? io_r_250_b : _GEN_13629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13631 = 9'hfb == r_count_33_io_out ? io_r_251_b : _GEN_13630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13632 = 9'hfc == r_count_33_io_out ? io_r_252_b : _GEN_13631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13633 = 9'hfd == r_count_33_io_out ? io_r_253_b : _GEN_13632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13634 = 9'hfe == r_count_33_io_out ? io_r_254_b : _GEN_13633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13635 = 9'hff == r_count_33_io_out ? io_r_255_b : _GEN_13634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13636 = 9'h100 == r_count_33_io_out ? io_r_256_b : _GEN_13635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13637 = 9'h101 == r_count_33_io_out ? io_r_257_b : _GEN_13636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13638 = 9'h102 == r_count_33_io_out ? io_r_258_b : _GEN_13637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13639 = 9'h103 == r_count_33_io_out ? io_r_259_b : _GEN_13638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13640 = 9'h104 == r_count_33_io_out ? io_r_260_b : _GEN_13639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13641 = 9'h105 == r_count_33_io_out ? io_r_261_b : _GEN_13640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13642 = 9'h106 == r_count_33_io_out ? io_r_262_b : _GEN_13641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13643 = 9'h107 == r_count_33_io_out ? io_r_263_b : _GEN_13642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13644 = 9'h108 == r_count_33_io_out ? io_r_264_b : _GEN_13643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13645 = 9'h109 == r_count_33_io_out ? io_r_265_b : _GEN_13644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13646 = 9'h10a == r_count_33_io_out ? io_r_266_b : _GEN_13645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13647 = 9'h10b == r_count_33_io_out ? io_r_267_b : _GEN_13646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13648 = 9'h10c == r_count_33_io_out ? io_r_268_b : _GEN_13647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13649 = 9'h10d == r_count_33_io_out ? io_r_269_b : _GEN_13648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13650 = 9'h10e == r_count_33_io_out ? io_r_270_b : _GEN_13649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13651 = 9'h10f == r_count_33_io_out ? io_r_271_b : _GEN_13650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13652 = 9'h110 == r_count_33_io_out ? io_r_272_b : _GEN_13651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13653 = 9'h111 == r_count_33_io_out ? io_r_273_b : _GEN_13652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13654 = 9'h112 == r_count_33_io_out ? io_r_274_b : _GEN_13653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13655 = 9'h113 == r_count_33_io_out ? io_r_275_b : _GEN_13654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13656 = 9'h114 == r_count_33_io_out ? io_r_276_b : _GEN_13655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13657 = 9'h115 == r_count_33_io_out ? io_r_277_b : _GEN_13656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13658 = 9'h116 == r_count_33_io_out ? io_r_278_b : _GEN_13657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13659 = 9'h117 == r_count_33_io_out ? io_r_279_b : _GEN_13658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13660 = 9'h118 == r_count_33_io_out ? io_r_280_b : _GEN_13659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13661 = 9'h119 == r_count_33_io_out ? io_r_281_b : _GEN_13660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13662 = 9'h11a == r_count_33_io_out ? io_r_282_b : _GEN_13661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13663 = 9'h11b == r_count_33_io_out ? io_r_283_b : _GEN_13662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13664 = 9'h11c == r_count_33_io_out ? io_r_284_b : _GEN_13663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13665 = 9'h11d == r_count_33_io_out ? io_r_285_b : _GEN_13664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13666 = 9'h11e == r_count_33_io_out ? io_r_286_b : _GEN_13665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13667 = 9'h11f == r_count_33_io_out ? io_r_287_b : _GEN_13666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13668 = 9'h120 == r_count_33_io_out ? io_r_288_b : _GEN_13667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13669 = 9'h121 == r_count_33_io_out ? io_r_289_b : _GEN_13668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13670 = 9'h122 == r_count_33_io_out ? io_r_290_b : _GEN_13669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13671 = 9'h123 == r_count_33_io_out ? io_r_291_b : _GEN_13670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13672 = 9'h124 == r_count_33_io_out ? io_r_292_b : _GEN_13671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13673 = 9'h125 == r_count_33_io_out ? io_r_293_b : _GEN_13672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13674 = 9'h126 == r_count_33_io_out ? io_r_294_b : _GEN_13673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13675 = 9'h127 == r_count_33_io_out ? io_r_295_b : _GEN_13674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13676 = 9'h128 == r_count_33_io_out ? io_r_296_b : _GEN_13675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13677 = 9'h129 == r_count_33_io_out ? io_r_297_b : _GEN_13676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13678 = 9'h12a == r_count_33_io_out ? io_r_298_b : _GEN_13677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13679 = 9'h12b == r_count_33_io_out ? io_r_299_b : _GEN_13678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13680 = 9'h12c == r_count_33_io_out ? io_r_300_b : _GEN_13679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13681 = 9'h12d == r_count_33_io_out ? io_r_301_b : _GEN_13680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13682 = 9'h12e == r_count_33_io_out ? io_r_302_b : _GEN_13681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13683 = 9'h12f == r_count_33_io_out ? io_r_303_b : _GEN_13682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13684 = 9'h130 == r_count_33_io_out ? io_r_304_b : _GEN_13683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13685 = 9'h131 == r_count_33_io_out ? io_r_305_b : _GEN_13684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13686 = 9'h132 == r_count_33_io_out ? io_r_306_b : _GEN_13685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13687 = 9'h133 == r_count_33_io_out ? io_r_307_b : _GEN_13686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13688 = 9'h134 == r_count_33_io_out ? io_r_308_b : _GEN_13687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13689 = 9'h135 == r_count_33_io_out ? io_r_309_b : _GEN_13688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13690 = 9'h136 == r_count_33_io_out ? io_r_310_b : _GEN_13689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13691 = 9'h137 == r_count_33_io_out ? io_r_311_b : _GEN_13690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13692 = 9'h138 == r_count_33_io_out ? io_r_312_b : _GEN_13691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13693 = 9'h139 == r_count_33_io_out ? io_r_313_b : _GEN_13692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13694 = 9'h13a == r_count_33_io_out ? io_r_314_b : _GEN_13693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13695 = 9'h13b == r_count_33_io_out ? io_r_315_b : _GEN_13694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13696 = 9'h13c == r_count_33_io_out ? io_r_316_b : _GEN_13695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13697 = 9'h13d == r_count_33_io_out ? io_r_317_b : _GEN_13696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13698 = 9'h13e == r_count_33_io_out ? io_r_318_b : _GEN_13697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13699 = 9'h13f == r_count_33_io_out ? io_r_319_b : _GEN_13698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13700 = 9'h140 == r_count_33_io_out ? io_r_320_b : _GEN_13699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13701 = 9'h141 == r_count_33_io_out ? io_r_321_b : _GEN_13700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13702 = 9'h142 == r_count_33_io_out ? io_r_322_b : _GEN_13701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13703 = 9'h143 == r_count_33_io_out ? io_r_323_b : _GEN_13702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13704 = 9'h144 == r_count_33_io_out ? io_r_324_b : _GEN_13703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13705 = 9'h145 == r_count_33_io_out ? io_r_325_b : _GEN_13704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13706 = 9'h146 == r_count_33_io_out ? io_r_326_b : _GEN_13705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13707 = 9'h147 == r_count_33_io_out ? io_r_327_b : _GEN_13706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13708 = 9'h148 == r_count_33_io_out ? io_r_328_b : _GEN_13707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13709 = 9'h149 == r_count_33_io_out ? io_r_329_b : _GEN_13708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13710 = 9'h14a == r_count_33_io_out ? io_r_330_b : _GEN_13709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13711 = 9'h14b == r_count_33_io_out ? io_r_331_b : _GEN_13710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13712 = 9'h14c == r_count_33_io_out ? io_r_332_b : _GEN_13711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13713 = 9'h14d == r_count_33_io_out ? io_r_333_b : _GEN_13712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13714 = 9'h14e == r_count_33_io_out ? io_r_334_b : _GEN_13713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13715 = 9'h14f == r_count_33_io_out ? io_r_335_b : _GEN_13714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13716 = 9'h150 == r_count_33_io_out ? io_r_336_b : _GEN_13715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13717 = 9'h151 == r_count_33_io_out ? io_r_337_b : _GEN_13716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13718 = 9'h152 == r_count_33_io_out ? io_r_338_b : _GEN_13717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13719 = 9'h153 == r_count_33_io_out ? io_r_339_b : _GEN_13718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13720 = 9'h154 == r_count_33_io_out ? io_r_340_b : _GEN_13719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13721 = 9'h155 == r_count_33_io_out ? io_r_341_b : _GEN_13720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13722 = 9'h156 == r_count_33_io_out ? io_r_342_b : _GEN_13721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13723 = 9'h157 == r_count_33_io_out ? io_r_343_b : _GEN_13722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13724 = 9'h158 == r_count_33_io_out ? io_r_344_b : _GEN_13723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13725 = 9'h159 == r_count_33_io_out ? io_r_345_b : _GEN_13724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13726 = 9'h15a == r_count_33_io_out ? io_r_346_b : _GEN_13725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13727 = 9'h15b == r_count_33_io_out ? io_r_347_b : _GEN_13726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13728 = 9'h15c == r_count_33_io_out ? io_r_348_b : _GEN_13727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13729 = 9'h15d == r_count_33_io_out ? io_r_349_b : _GEN_13728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13730 = 9'h15e == r_count_33_io_out ? io_r_350_b : _GEN_13729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13731 = 9'h15f == r_count_33_io_out ? io_r_351_b : _GEN_13730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13732 = 9'h160 == r_count_33_io_out ? io_r_352_b : _GEN_13731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13733 = 9'h161 == r_count_33_io_out ? io_r_353_b : _GEN_13732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13734 = 9'h162 == r_count_33_io_out ? io_r_354_b : _GEN_13733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13735 = 9'h163 == r_count_33_io_out ? io_r_355_b : _GEN_13734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13736 = 9'h164 == r_count_33_io_out ? io_r_356_b : _GEN_13735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13737 = 9'h165 == r_count_33_io_out ? io_r_357_b : _GEN_13736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13738 = 9'h166 == r_count_33_io_out ? io_r_358_b : _GEN_13737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13739 = 9'h167 == r_count_33_io_out ? io_r_359_b : _GEN_13738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13740 = 9'h168 == r_count_33_io_out ? io_r_360_b : _GEN_13739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13741 = 9'h169 == r_count_33_io_out ? io_r_361_b : _GEN_13740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13742 = 9'h16a == r_count_33_io_out ? io_r_362_b : _GEN_13741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13743 = 9'h16b == r_count_33_io_out ? io_r_363_b : _GEN_13742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13744 = 9'h16c == r_count_33_io_out ? io_r_364_b : _GEN_13743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13745 = 9'h16d == r_count_33_io_out ? io_r_365_b : _GEN_13744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13746 = 9'h16e == r_count_33_io_out ? io_r_366_b : _GEN_13745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13747 = 9'h16f == r_count_33_io_out ? io_r_367_b : _GEN_13746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13748 = 9'h170 == r_count_33_io_out ? io_r_368_b : _GEN_13747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13749 = 9'h171 == r_count_33_io_out ? io_r_369_b : _GEN_13748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13750 = 9'h172 == r_count_33_io_out ? io_r_370_b : _GEN_13749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13751 = 9'h173 == r_count_33_io_out ? io_r_371_b : _GEN_13750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13752 = 9'h174 == r_count_33_io_out ? io_r_372_b : _GEN_13751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13753 = 9'h175 == r_count_33_io_out ? io_r_373_b : _GEN_13752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13754 = 9'h176 == r_count_33_io_out ? io_r_374_b : _GEN_13753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13755 = 9'h177 == r_count_33_io_out ? io_r_375_b : _GEN_13754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13756 = 9'h178 == r_count_33_io_out ? io_r_376_b : _GEN_13755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13757 = 9'h179 == r_count_33_io_out ? io_r_377_b : _GEN_13756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13758 = 9'h17a == r_count_33_io_out ? io_r_378_b : _GEN_13757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13759 = 9'h17b == r_count_33_io_out ? io_r_379_b : _GEN_13758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13760 = 9'h17c == r_count_33_io_out ? io_r_380_b : _GEN_13759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13761 = 9'h17d == r_count_33_io_out ? io_r_381_b : _GEN_13760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13762 = 9'h17e == r_count_33_io_out ? io_r_382_b : _GEN_13761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13763 = 9'h17f == r_count_33_io_out ? io_r_383_b : _GEN_13762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13764 = 9'h180 == r_count_33_io_out ? io_r_384_b : _GEN_13763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13765 = 9'h181 == r_count_33_io_out ? io_r_385_b : _GEN_13764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13766 = 9'h182 == r_count_33_io_out ? io_r_386_b : _GEN_13765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13767 = 9'h183 == r_count_33_io_out ? io_r_387_b : _GEN_13766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13768 = 9'h184 == r_count_33_io_out ? io_r_388_b : _GEN_13767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13769 = 9'h185 == r_count_33_io_out ? io_r_389_b : _GEN_13768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13770 = 9'h186 == r_count_33_io_out ? io_r_390_b : _GEN_13769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13771 = 9'h187 == r_count_33_io_out ? io_r_391_b : _GEN_13770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13772 = 9'h188 == r_count_33_io_out ? io_r_392_b : _GEN_13771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13773 = 9'h189 == r_count_33_io_out ? io_r_393_b : _GEN_13772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13774 = 9'h18a == r_count_33_io_out ? io_r_394_b : _GEN_13773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13775 = 9'h18b == r_count_33_io_out ? io_r_395_b : _GEN_13774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13776 = 9'h18c == r_count_33_io_out ? io_r_396_b : _GEN_13775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13777 = 9'h18d == r_count_33_io_out ? io_r_397_b : _GEN_13776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13778 = 9'h18e == r_count_33_io_out ? io_r_398_b : _GEN_13777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13781 = 9'h1 == r_count_34_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13782 = 9'h2 == r_count_34_io_out ? io_r_2_b : _GEN_13781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13783 = 9'h3 == r_count_34_io_out ? io_r_3_b : _GEN_13782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13784 = 9'h4 == r_count_34_io_out ? io_r_4_b : _GEN_13783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13785 = 9'h5 == r_count_34_io_out ? io_r_5_b : _GEN_13784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13786 = 9'h6 == r_count_34_io_out ? io_r_6_b : _GEN_13785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13787 = 9'h7 == r_count_34_io_out ? io_r_7_b : _GEN_13786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13788 = 9'h8 == r_count_34_io_out ? io_r_8_b : _GEN_13787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13789 = 9'h9 == r_count_34_io_out ? io_r_9_b : _GEN_13788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13790 = 9'ha == r_count_34_io_out ? io_r_10_b : _GEN_13789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13791 = 9'hb == r_count_34_io_out ? io_r_11_b : _GEN_13790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13792 = 9'hc == r_count_34_io_out ? io_r_12_b : _GEN_13791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13793 = 9'hd == r_count_34_io_out ? io_r_13_b : _GEN_13792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13794 = 9'he == r_count_34_io_out ? io_r_14_b : _GEN_13793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13795 = 9'hf == r_count_34_io_out ? io_r_15_b : _GEN_13794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13796 = 9'h10 == r_count_34_io_out ? io_r_16_b : _GEN_13795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13797 = 9'h11 == r_count_34_io_out ? io_r_17_b : _GEN_13796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13798 = 9'h12 == r_count_34_io_out ? io_r_18_b : _GEN_13797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13799 = 9'h13 == r_count_34_io_out ? io_r_19_b : _GEN_13798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13800 = 9'h14 == r_count_34_io_out ? io_r_20_b : _GEN_13799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13801 = 9'h15 == r_count_34_io_out ? io_r_21_b : _GEN_13800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13802 = 9'h16 == r_count_34_io_out ? io_r_22_b : _GEN_13801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13803 = 9'h17 == r_count_34_io_out ? io_r_23_b : _GEN_13802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13804 = 9'h18 == r_count_34_io_out ? io_r_24_b : _GEN_13803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13805 = 9'h19 == r_count_34_io_out ? io_r_25_b : _GEN_13804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13806 = 9'h1a == r_count_34_io_out ? io_r_26_b : _GEN_13805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13807 = 9'h1b == r_count_34_io_out ? io_r_27_b : _GEN_13806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13808 = 9'h1c == r_count_34_io_out ? io_r_28_b : _GEN_13807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13809 = 9'h1d == r_count_34_io_out ? io_r_29_b : _GEN_13808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13810 = 9'h1e == r_count_34_io_out ? io_r_30_b : _GEN_13809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13811 = 9'h1f == r_count_34_io_out ? io_r_31_b : _GEN_13810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13812 = 9'h20 == r_count_34_io_out ? io_r_32_b : _GEN_13811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13813 = 9'h21 == r_count_34_io_out ? io_r_33_b : _GEN_13812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13814 = 9'h22 == r_count_34_io_out ? io_r_34_b : _GEN_13813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13815 = 9'h23 == r_count_34_io_out ? io_r_35_b : _GEN_13814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13816 = 9'h24 == r_count_34_io_out ? io_r_36_b : _GEN_13815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13817 = 9'h25 == r_count_34_io_out ? io_r_37_b : _GEN_13816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13818 = 9'h26 == r_count_34_io_out ? io_r_38_b : _GEN_13817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13819 = 9'h27 == r_count_34_io_out ? io_r_39_b : _GEN_13818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13820 = 9'h28 == r_count_34_io_out ? io_r_40_b : _GEN_13819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13821 = 9'h29 == r_count_34_io_out ? io_r_41_b : _GEN_13820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13822 = 9'h2a == r_count_34_io_out ? io_r_42_b : _GEN_13821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13823 = 9'h2b == r_count_34_io_out ? io_r_43_b : _GEN_13822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13824 = 9'h2c == r_count_34_io_out ? io_r_44_b : _GEN_13823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13825 = 9'h2d == r_count_34_io_out ? io_r_45_b : _GEN_13824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13826 = 9'h2e == r_count_34_io_out ? io_r_46_b : _GEN_13825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13827 = 9'h2f == r_count_34_io_out ? io_r_47_b : _GEN_13826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13828 = 9'h30 == r_count_34_io_out ? io_r_48_b : _GEN_13827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13829 = 9'h31 == r_count_34_io_out ? io_r_49_b : _GEN_13828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13830 = 9'h32 == r_count_34_io_out ? io_r_50_b : _GEN_13829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13831 = 9'h33 == r_count_34_io_out ? io_r_51_b : _GEN_13830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13832 = 9'h34 == r_count_34_io_out ? io_r_52_b : _GEN_13831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13833 = 9'h35 == r_count_34_io_out ? io_r_53_b : _GEN_13832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13834 = 9'h36 == r_count_34_io_out ? io_r_54_b : _GEN_13833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13835 = 9'h37 == r_count_34_io_out ? io_r_55_b : _GEN_13834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13836 = 9'h38 == r_count_34_io_out ? io_r_56_b : _GEN_13835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13837 = 9'h39 == r_count_34_io_out ? io_r_57_b : _GEN_13836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13838 = 9'h3a == r_count_34_io_out ? io_r_58_b : _GEN_13837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13839 = 9'h3b == r_count_34_io_out ? io_r_59_b : _GEN_13838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13840 = 9'h3c == r_count_34_io_out ? io_r_60_b : _GEN_13839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13841 = 9'h3d == r_count_34_io_out ? io_r_61_b : _GEN_13840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13842 = 9'h3e == r_count_34_io_out ? io_r_62_b : _GEN_13841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13843 = 9'h3f == r_count_34_io_out ? io_r_63_b : _GEN_13842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13844 = 9'h40 == r_count_34_io_out ? io_r_64_b : _GEN_13843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13845 = 9'h41 == r_count_34_io_out ? io_r_65_b : _GEN_13844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13846 = 9'h42 == r_count_34_io_out ? io_r_66_b : _GEN_13845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13847 = 9'h43 == r_count_34_io_out ? io_r_67_b : _GEN_13846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13848 = 9'h44 == r_count_34_io_out ? io_r_68_b : _GEN_13847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13849 = 9'h45 == r_count_34_io_out ? io_r_69_b : _GEN_13848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13850 = 9'h46 == r_count_34_io_out ? io_r_70_b : _GEN_13849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13851 = 9'h47 == r_count_34_io_out ? io_r_71_b : _GEN_13850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13852 = 9'h48 == r_count_34_io_out ? io_r_72_b : _GEN_13851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13853 = 9'h49 == r_count_34_io_out ? io_r_73_b : _GEN_13852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13854 = 9'h4a == r_count_34_io_out ? io_r_74_b : _GEN_13853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13855 = 9'h4b == r_count_34_io_out ? io_r_75_b : _GEN_13854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13856 = 9'h4c == r_count_34_io_out ? io_r_76_b : _GEN_13855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13857 = 9'h4d == r_count_34_io_out ? io_r_77_b : _GEN_13856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13858 = 9'h4e == r_count_34_io_out ? io_r_78_b : _GEN_13857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13859 = 9'h4f == r_count_34_io_out ? io_r_79_b : _GEN_13858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13860 = 9'h50 == r_count_34_io_out ? io_r_80_b : _GEN_13859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13861 = 9'h51 == r_count_34_io_out ? io_r_81_b : _GEN_13860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13862 = 9'h52 == r_count_34_io_out ? io_r_82_b : _GEN_13861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13863 = 9'h53 == r_count_34_io_out ? io_r_83_b : _GEN_13862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13864 = 9'h54 == r_count_34_io_out ? io_r_84_b : _GEN_13863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13865 = 9'h55 == r_count_34_io_out ? io_r_85_b : _GEN_13864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13866 = 9'h56 == r_count_34_io_out ? io_r_86_b : _GEN_13865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13867 = 9'h57 == r_count_34_io_out ? io_r_87_b : _GEN_13866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13868 = 9'h58 == r_count_34_io_out ? io_r_88_b : _GEN_13867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13869 = 9'h59 == r_count_34_io_out ? io_r_89_b : _GEN_13868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13870 = 9'h5a == r_count_34_io_out ? io_r_90_b : _GEN_13869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13871 = 9'h5b == r_count_34_io_out ? io_r_91_b : _GEN_13870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13872 = 9'h5c == r_count_34_io_out ? io_r_92_b : _GEN_13871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13873 = 9'h5d == r_count_34_io_out ? io_r_93_b : _GEN_13872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13874 = 9'h5e == r_count_34_io_out ? io_r_94_b : _GEN_13873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13875 = 9'h5f == r_count_34_io_out ? io_r_95_b : _GEN_13874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13876 = 9'h60 == r_count_34_io_out ? io_r_96_b : _GEN_13875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13877 = 9'h61 == r_count_34_io_out ? io_r_97_b : _GEN_13876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13878 = 9'h62 == r_count_34_io_out ? io_r_98_b : _GEN_13877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13879 = 9'h63 == r_count_34_io_out ? io_r_99_b : _GEN_13878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13880 = 9'h64 == r_count_34_io_out ? io_r_100_b : _GEN_13879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13881 = 9'h65 == r_count_34_io_out ? io_r_101_b : _GEN_13880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13882 = 9'h66 == r_count_34_io_out ? io_r_102_b : _GEN_13881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13883 = 9'h67 == r_count_34_io_out ? io_r_103_b : _GEN_13882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13884 = 9'h68 == r_count_34_io_out ? io_r_104_b : _GEN_13883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13885 = 9'h69 == r_count_34_io_out ? io_r_105_b : _GEN_13884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13886 = 9'h6a == r_count_34_io_out ? io_r_106_b : _GEN_13885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13887 = 9'h6b == r_count_34_io_out ? io_r_107_b : _GEN_13886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13888 = 9'h6c == r_count_34_io_out ? io_r_108_b : _GEN_13887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13889 = 9'h6d == r_count_34_io_out ? io_r_109_b : _GEN_13888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13890 = 9'h6e == r_count_34_io_out ? io_r_110_b : _GEN_13889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13891 = 9'h6f == r_count_34_io_out ? io_r_111_b : _GEN_13890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13892 = 9'h70 == r_count_34_io_out ? io_r_112_b : _GEN_13891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13893 = 9'h71 == r_count_34_io_out ? io_r_113_b : _GEN_13892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13894 = 9'h72 == r_count_34_io_out ? io_r_114_b : _GEN_13893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13895 = 9'h73 == r_count_34_io_out ? io_r_115_b : _GEN_13894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13896 = 9'h74 == r_count_34_io_out ? io_r_116_b : _GEN_13895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13897 = 9'h75 == r_count_34_io_out ? io_r_117_b : _GEN_13896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13898 = 9'h76 == r_count_34_io_out ? io_r_118_b : _GEN_13897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13899 = 9'h77 == r_count_34_io_out ? io_r_119_b : _GEN_13898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13900 = 9'h78 == r_count_34_io_out ? io_r_120_b : _GEN_13899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13901 = 9'h79 == r_count_34_io_out ? io_r_121_b : _GEN_13900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13902 = 9'h7a == r_count_34_io_out ? io_r_122_b : _GEN_13901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13903 = 9'h7b == r_count_34_io_out ? io_r_123_b : _GEN_13902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13904 = 9'h7c == r_count_34_io_out ? io_r_124_b : _GEN_13903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13905 = 9'h7d == r_count_34_io_out ? io_r_125_b : _GEN_13904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13906 = 9'h7e == r_count_34_io_out ? io_r_126_b : _GEN_13905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13907 = 9'h7f == r_count_34_io_out ? io_r_127_b : _GEN_13906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13908 = 9'h80 == r_count_34_io_out ? io_r_128_b : _GEN_13907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13909 = 9'h81 == r_count_34_io_out ? io_r_129_b : _GEN_13908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13910 = 9'h82 == r_count_34_io_out ? io_r_130_b : _GEN_13909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13911 = 9'h83 == r_count_34_io_out ? io_r_131_b : _GEN_13910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13912 = 9'h84 == r_count_34_io_out ? io_r_132_b : _GEN_13911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13913 = 9'h85 == r_count_34_io_out ? io_r_133_b : _GEN_13912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13914 = 9'h86 == r_count_34_io_out ? io_r_134_b : _GEN_13913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13915 = 9'h87 == r_count_34_io_out ? io_r_135_b : _GEN_13914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13916 = 9'h88 == r_count_34_io_out ? io_r_136_b : _GEN_13915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13917 = 9'h89 == r_count_34_io_out ? io_r_137_b : _GEN_13916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13918 = 9'h8a == r_count_34_io_out ? io_r_138_b : _GEN_13917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13919 = 9'h8b == r_count_34_io_out ? io_r_139_b : _GEN_13918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13920 = 9'h8c == r_count_34_io_out ? io_r_140_b : _GEN_13919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13921 = 9'h8d == r_count_34_io_out ? io_r_141_b : _GEN_13920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13922 = 9'h8e == r_count_34_io_out ? io_r_142_b : _GEN_13921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13923 = 9'h8f == r_count_34_io_out ? io_r_143_b : _GEN_13922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13924 = 9'h90 == r_count_34_io_out ? io_r_144_b : _GEN_13923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13925 = 9'h91 == r_count_34_io_out ? io_r_145_b : _GEN_13924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13926 = 9'h92 == r_count_34_io_out ? io_r_146_b : _GEN_13925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13927 = 9'h93 == r_count_34_io_out ? io_r_147_b : _GEN_13926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13928 = 9'h94 == r_count_34_io_out ? io_r_148_b : _GEN_13927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13929 = 9'h95 == r_count_34_io_out ? io_r_149_b : _GEN_13928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13930 = 9'h96 == r_count_34_io_out ? io_r_150_b : _GEN_13929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13931 = 9'h97 == r_count_34_io_out ? io_r_151_b : _GEN_13930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13932 = 9'h98 == r_count_34_io_out ? io_r_152_b : _GEN_13931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13933 = 9'h99 == r_count_34_io_out ? io_r_153_b : _GEN_13932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13934 = 9'h9a == r_count_34_io_out ? io_r_154_b : _GEN_13933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13935 = 9'h9b == r_count_34_io_out ? io_r_155_b : _GEN_13934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13936 = 9'h9c == r_count_34_io_out ? io_r_156_b : _GEN_13935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13937 = 9'h9d == r_count_34_io_out ? io_r_157_b : _GEN_13936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13938 = 9'h9e == r_count_34_io_out ? io_r_158_b : _GEN_13937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13939 = 9'h9f == r_count_34_io_out ? io_r_159_b : _GEN_13938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13940 = 9'ha0 == r_count_34_io_out ? io_r_160_b : _GEN_13939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13941 = 9'ha1 == r_count_34_io_out ? io_r_161_b : _GEN_13940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13942 = 9'ha2 == r_count_34_io_out ? io_r_162_b : _GEN_13941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13943 = 9'ha3 == r_count_34_io_out ? io_r_163_b : _GEN_13942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13944 = 9'ha4 == r_count_34_io_out ? io_r_164_b : _GEN_13943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13945 = 9'ha5 == r_count_34_io_out ? io_r_165_b : _GEN_13944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13946 = 9'ha6 == r_count_34_io_out ? io_r_166_b : _GEN_13945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13947 = 9'ha7 == r_count_34_io_out ? io_r_167_b : _GEN_13946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13948 = 9'ha8 == r_count_34_io_out ? io_r_168_b : _GEN_13947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13949 = 9'ha9 == r_count_34_io_out ? io_r_169_b : _GEN_13948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13950 = 9'haa == r_count_34_io_out ? io_r_170_b : _GEN_13949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13951 = 9'hab == r_count_34_io_out ? io_r_171_b : _GEN_13950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13952 = 9'hac == r_count_34_io_out ? io_r_172_b : _GEN_13951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13953 = 9'had == r_count_34_io_out ? io_r_173_b : _GEN_13952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13954 = 9'hae == r_count_34_io_out ? io_r_174_b : _GEN_13953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13955 = 9'haf == r_count_34_io_out ? io_r_175_b : _GEN_13954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13956 = 9'hb0 == r_count_34_io_out ? io_r_176_b : _GEN_13955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13957 = 9'hb1 == r_count_34_io_out ? io_r_177_b : _GEN_13956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13958 = 9'hb2 == r_count_34_io_out ? io_r_178_b : _GEN_13957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13959 = 9'hb3 == r_count_34_io_out ? io_r_179_b : _GEN_13958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13960 = 9'hb4 == r_count_34_io_out ? io_r_180_b : _GEN_13959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13961 = 9'hb5 == r_count_34_io_out ? io_r_181_b : _GEN_13960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13962 = 9'hb6 == r_count_34_io_out ? io_r_182_b : _GEN_13961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13963 = 9'hb7 == r_count_34_io_out ? io_r_183_b : _GEN_13962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13964 = 9'hb8 == r_count_34_io_out ? io_r_184_b : _GEN_13963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13965 = 9'hb9 == r_count_34_io_out ? io_r_185_b : _GEN_13964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13966 = 9'hba == r_count_34_io_out ? io_r_186_b : _GEN_13965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13967 = 9'hbb == r_count_34_io_out ? io_r_187_b : _GEN_13966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13968 = 9'hbc == r_count_34_io_out ? io_r_188_b : _GEN_13967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13969 = 9'hbd == r_count_34_io_out ? io_r_189_b : _GEN_13968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13970 = 9'hbe == r_count_34_io_out ? io_r_190_b : _GEN_13969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13971 = 9'hbf == r_count_34_io_out ? io_r_191_b : _GEN_13970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13972 = 9'hc0 == r_count_34_io_out ? io_r_192_b : _GEN_13971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13973 = 9'hc1 == r_count_34_io_out ? io_r_193_b : _GEN_13972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13974 = 9'hc2 == r_count_34_io_out ? io_r_194_b : _GEN_13973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13975 = 9'hc3 == r_count_34_io_out ? io_r_195_b : _GEN_13974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13976 = 9'hc4 == r_count_34_io_out ? io_r_196_b : _GEN_13975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13977 = 9'hc5 == r_count_34_io_out ? io_r_197_b : _GEN_13976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13978 = 9'hc6 == r_count_34_io_out ? io_r_198_b : _GEN_13977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13979 = 9'hc7 == r_count_34_io_out ? io_r_199_b : _GEN_13978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13980 = 9'hc8 == r_count_34_io_out ? io_r_200_b : _GEN_13979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13981 = 9'hc9 == r_count_34_io_out ? io_r_201_b : _GEN_13980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13982 = 9'hca == r_count_34_io_out ? io_r_202_b : _GEN_13981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13983 = 9'hcb == r_count_34_io_out ? io_r_203_b : _GEN_13982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13984 = 9'hcc == r_count_34_io_out ? io_r_204_b : _GEN_13983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13985 = 9'hcd == r_count_34_io_out ? io_r_205_b : _GEN_13984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13986 = 9'hce == r_count_34_io_out ? io_r_206_b : _GEN_13985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13987 = 9'hcf == r_count_34_io_out ? io_r_207_b : _GEN_13986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13988 = 9'hd0 == r_count_34_io_out ? io_r_208_b : _GEN_13987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13989 = 9'hd1 == r_count_34_io_out ? io_r_209_b : _GEN_13988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13990 = 9'hd2 == r_count_34_io_out ? io_r_210_b : _GEN_13989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13991 = 9'hd3 == r_count_34_io_out ? io_r_211_b : _GEN_13990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13992 = 9'hd4 == r_count_34_io_out ? io_r_212_b : _GEN_13991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13993 = 9'hd5 == r_count_34_io_out ? io_r_213_b : _GEN_13992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13994 = 9'hd6 == r_count_34_io_out ? io_r_214_b : _GEN_13993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13995 = 9'hd7 == r_count_34_io_out ? io_r_215_b : _GEN_13994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13996 = 9'hd8 == r_count_34_io_out ? io_r_216_b : _GEN_13995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13997 = 9'hd9 == r_count_34_io_out ? io_r_217_b : _GEN_13996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13998 = 9'hda == r_count_34_io_out ? io_r_218_b : _GEN_13997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13999 = 9'hdb == r_count_34_io_out ? io_r_219_b : _GEN_13998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14000 = 9'hdc == r_count_34_io_out ? io_r_220_b : _GEN_13999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14001 = 9'hdd == r_count_34_io_out ? io_r_221_b : _GEN_14000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14002 = 9'hde == r_count_34_io_out ? io_r_222_b : _GEN_14001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14003 = 9'hdf == r_count_34_io_out ? io_r_223_b : _GEN_14002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14004 = 9'he0 == r_count_34_io_out ? io_r_224_b : _GEN_14003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14005 = 9'he1 == r_count_34_io_out ? io_r_225_b : _GEN_14004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14006 = 9'he2 == r_count_34_io_out ? io_r_226_b : _GEN_14005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14007 = 9'he3 == r_count_34_io_out ? io_r_227_b : _GEN_14006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14008 = 9'he4 == r_count_34_io_out ? io_r_228_b : _GEN_14007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14009 = 9'he5 == r_count_34_io_out ? io_r_229_b : _GEN_14008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14010 = 9'he6 == r_count_34_io_out ? io_r_230_b : _GEN_14009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14011 = 9'he7 == r_count_34_io_out ? io_r_231_b : _GEN_14010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14012 = 9'he8 == r_count_34_io_out ? io_r_232_b : _GEN_14011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14013 = 9'he9 == r_count_34_io_out ? io_r_233_b : _GEN_14012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14014 = 9'hea == r_count_34_io_out ? io_r_234_b : _GEN_14013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14015 = 9'heb == r_count_34_io_out ? io_r_235_b : _GEN_14014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14016 = 9'hec == r_count_34_io_out ? io_r_236_b : _GEN_14015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14017 = 9'hed == r_count_34_io_out ? io_r_237_b : _GEN_14016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14018 = 9'hee == r_count_34_io_out ? io_r_238_b : _GEN_14017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14019 = 9'hef == r_count_34_io_out ? io_r_239_b : _GEN_14018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14020 = 9'hf0 == r_count_34_io_out ? io_r_240_b : _GEN_14019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14021 = 9'hf1 == r_count_34_io_out ? io_r_241_b : _GEN_14020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14022 = 9'hf2 == r_count_34_io_out ? io_r_242_b : _GEN_14021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14023 = 9'hf3 == r_count_34_io_out ? io_r_243_b : _GEN_14022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14024 = 9'hf4 == r_count_34_io_out ? io_r_244_b : _GEN_14023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14025 = 9'hf5 == r_count_34_io_out ? io_r_245_b : _GEN_14024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14026 = 9'hf6 == r_count_34_io_out ? io_r_246_b : _GEN_14025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14027 = 9'hf7 == r_count_34_io_out ? io_r_247_b : _GEN_14026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14028 = 9'hf8 == r_count_34_io_out ? io_r_248_b : _GEN_14027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14029 = 9'hf9 == r_count_34_io_out ? io_r_249_b : _GEN_14028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14030 = 9'hfa == r_count_34_io_out ? io_r_250_b : _GEN_14029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14031 = 9'hfb == r_count_34_io_out ? io_r_251_b : _GEN_14030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14032 = 9'hfc == r_count_34_io_out ? io_r_252_b : _GEN_14031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14033 = 9'hfd == r_count_34_io_out ? io_r_253_b : _GEN_14032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14034 = 9'hfe == r_count_34_io_out ? io_r_254_b : _GEN_14033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14035 = 9'hff == r_count_34_io_out ? io_r_255_b : _GEN_14034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14036 = 9'h100 == r_count_34_io_out ? io_r_256_b : _GEN_14035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14037 = 9'h101 == r_count_34_io_out ? io_r_257_b : _GEN_14036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14038 = 9'h102 == r_count_34_io_out ? io_r_258_b : _GEN_14037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14039 = 9'h103 == r_count_34_io_out ? io_r_259_b : _GEN_14038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14040 = 9'h104 == r_count_34_io_out ? io_r_260_b : _GEN_14039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14041 = 9'h105 == r_count_34_io_out ? io_r_261_b : _GEN_14040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14042 = 9'h106 == r_count_34_io_out ? io_r_262_b : _GEN_14041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14043 = 9'h107 == r_count_34_io_out ? io_r_263_b : _GEN_14042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14044 = 9'h108 == r_count_34_io_out ? io_r_264_b : _GEN_14043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14045 = 9'h109 == r_count_34_io_out ? io_r_265_b : _GEN_14044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14046 = 9'h10a == r_count_34_io_out ? io_r_266_b : _GEN_14045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14047 = 9'h10b == r_count_34_io_out ? io_r_267_b : _GEN_14046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14048 = 9'h10c == r_count_34_io_out ? io_r_268_b : _GEN_14047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14049 = 9'h10d == r_count_34_io_out ? io_r_269_b : _GEN_14048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14050 = 9'h10e == r_count_34_io_out ? io_r_270_b : _GEN_14049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14051 = 9'h10f == r_count_34_io_out ? io_r_271_b : _GEN_14050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14052 = 9'h110 == r_count_34_io_out ? io_r_272_b : _GEN_14051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14053 = 9'h111 == r_count_34_io_out ? io_r_273_b : _GEN_14052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14054 = 9'h112 == r_count_34_io_out ? io_r_274_b : _GEN_14053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14055 = 9'h113 == r_count_34_io_out ? io_r_275_b : _GEN_14054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14056 = 9'h114 == r_count_34_io_out ? io_r_276_b : _GEN_14055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14057 = 9'h115 == r_count_34_io_out ? io_r_277_b : _GEN_14056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14058 = 9'h116 == r_count_34_io_out ? io_r_278_b : _GEN_14057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14059 = 9'h117 == r_count_34_io_out ? io_r_279_b : _GEN_14058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14060 = 9'h118 == r_count_34_io_out ? io_r_280_b : _GEN_14059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14061 = 9'h119 == r_count_34_io_out ? io_r_281_b : _GEN_14060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14062 = 9'h11a == r_count_34_io_out ? io_r_282_b : _GEN_14061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14063 = 9'h11b == r_count_34_io_out ? io_r_283_b : _GEN_14062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14064 = 9'h11c == r_count_34_io_out ? io_r_284_b : _GEN_14063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14065 = 9'h11d == r_count_34_io_out ? io_r_285_b : _GEN_14064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14066 = 9'h11e == r_count_34_io_out ? io_r_286_b : _GEN_14065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14067 = 9'h11f == r_count_34_io_out ? io_r_287_b : _GEN_14066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14068 = 9'h120 == r_count_34_io_out ? io_r_288_b : _GEN_14067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14069 = 9'h121 == r_count_34_io_out ? io_r_289_b : _GEN_14068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14070 = 9'h122 == r_count_34_io_out ? io_r_290_b : _GEN_14069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14071 = 9'h123 == r_count_34_io_out ? io_r_291_b : _GEN_14070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14072 = 9'h124 == r_count_34_io_out ? io_r_292_b : _GEN_14071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14073 = 9'h125 == r_count_34_io_out ? io_r_293_b : _GEN_14072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14074 = 9'h126 == r_count_34_io_out ? io_r_294_b : _GEN_14073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14075 = 9'h127 == r_count_34_io_out ? io_r_295_b : _GEN_14074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14076 = 9'h128 == r_count_34_io_out ? io_r_296_b : _GEN_14075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14077 = 9'h129 == r_count_34_io_out ? io_r_297_b : _GEN_14076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14078 = 9'h12a == r_count_34_io_out ? io_r_298_b : _GEN_14077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14079 = 9'h12b == r_count_34_io_out ? io_r_299_b : _GEN_14078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14080 = 9'h12c == r_count_34_io_out ? io_r_300_b : _GEN_14079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14081 = 9'h12d == r_count_34_io_out ? io_r_301_b : _GEN_14080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14082 = 9'h12e == r_count_34_io_out ? io_r_302_b : _GEN_14081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14083 = 9'h12f == r_count_34_io_out ? io_r_303_b : _GEN_14082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14084 = 9'h130 == r_count_34_io_out ? io_r_304_b : _GEN_14083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14085 = 9'h131 == r_count_34_io_out ? io_r_305_b : _GEN_14084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14086 = 9'h132 == r_count_34_io_out ? io_r_306_b : _GEN_14085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14087 = 9'h133 == r_count_34_io_out ? io_r_307_b : _GEN_14086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14088 = 9'h134 == r_count_34_io_out ? io_r_308_b : _GEN_14087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14089 = 9'h135 == r_count_34_io_out ? io_r_309_b : _GEN_14088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14090 = 9'h136 == r_count_34_io_out ? io_r_310_b : _GEN_14089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14091 = 9'h137 == r_count_34_io_out ? io_r_311_b : _GEN_14090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14092 = 9'h138 == r_count_34_io_out ? io_r_312_b : _GEN_14091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14093 = 9'h139 == r_count_34_io_out ? io_r_313_b : _GEN_14092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14094 = 9'h13a == r_count_34_io_out ? io_r_314_b : _GEN_14093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14095 = 9'h13b == r_count_34_io_out ? io_r_315_b : _GEN_14094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14096 = 9'h13c == r_count_34_io_out ? io_r_316_b : _GEN_14095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14097 = 9'h13d == r_count_34_io_out ? io_r_317_b : _GEN_14096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14098 = 9'h13e == r_count_34_io_out ? io_r_318_b : _GEN_14097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14099 = 9'h13f == r_count_34_io_out ? io_r_319_b : _GEN_14098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14100 = 9'h140 == r_count_34_io_out ? io_r_320_b : _GEN_14099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14101 = 9'h141 == r_count_34_io_out ? io_r_321_b : _GEN_14100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14102 = 9'h142 == r_count_34_io_out ? io_r_322_b : _GEN_14101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14103 = 9'h143 == r_count_34_io_out ? io_r_323_b : _GEN_14102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14104 = 9'h144 == r_count_34_io_out ? io_r_324_b : _GEN_14103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14105 = 9'h145 == r_count_34_io_out ? io_r_325_b : _GEN_14104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14106 = 9'h146 == r_count_34_io_out ? io_r_326_b : _GEN_14105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14107 = 9'h147 == r_count_34_io_out ? io_r_327_b : _GEN_14106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14108 = 9'h148 == r_count_34_io_out ? io_r_328_b : _GEN_14107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14109 = 9'h149 == r_count_34_io_out ? io_r_329_b : _GEN_14108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14110 = 9'h14a == r_count_34_io_out ? io_r_330_b : _GEN_14109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14111 = 9'h14b == r_count_34_io_out ? io_r_331_b : _GEN_14110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14112 = 9'h14c == r_count_34_io_out ? io_r_332_b : _GEN_14111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14113 = 9'h14d == r_count_34_io_out ? io_r_333_b : _GEN_14112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14114 = 9'h14e == r_count_34_io_out ? io_r_334_b : _GEN_14113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14115 = 9'h14f == r_count_34_io_out ? io_r_335_b : _GEN_14114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14116 = 9'h150 == r_count_34_io_out ? io_r_336_b : _GEN_14115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14117 = 9'h151 == r_count_34_io_out ? io_r_337_b : _GEN_14116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14118 = 9'h152 == r_count_34_io_out ? io_r_338_b : _GEN_14117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14119 = 9'h153 == r_count_34_io_out ? io_r_339_b : _GEN_14118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14120 = 9'h154 == r_count_34_io_out ? io_r_340_b : _GEN_14119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14121 = 9'h155 == r_count_34_io_out ? io_r_341_b : _GEN_14120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14122 = 9'h156 == r_count_34_io_out ? io_r_342_b : _GEN_14121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14123 = 9'h157 == r_count_34_io_out ? io_r_343_b : _GEN_14122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14124 = 9'h158 == r_count_34_io_out ? io_r_344_b : _GEN_14123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14125 = 9'h159 == r_count_34_io_out ? io_r_345_b : _GEN_14124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14126 = 9'h15a == r_count_34_io_out ? io_r_346_b : _GEN_14125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14127 = 9'h15b == r_count_34_io_out ? io_r_347_b : _GEN_14126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14128 = 9'h15c == r_count_34_io_out ? io_r_348_b : _GEN_14127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14129 = 9'h15d == r_count_34_io_out ? io_r_349_b : _GEN_14128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14130 = 9'h15e == r_count_34_io_out ? io_r_350_b : _GEN_14129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14131 = 9'h15f == r_count_34_io_out ? io_r_351_b : _GEN_14130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14132 = 9'h160 == r_count_34_io_out ? io_r_352_b : _GEN_14131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14133 = 9'h161 == r_count_34_io_out ? io_r_353_b : _GEN_14132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14134 = 9'h162 == r_count_34_io_out ? io_r_354_b : _GEN_14133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14135 = 9'h163 == r_count_34_io_out ? io_r_355_b : _GEN_14134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14136 = 9'h164 == r_count_34_io_out ? io_r_356_b : _GEN_14135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14137 = 9'h165 == r_count_34_io_out ? io_r_357_b : _GEN_14136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14138 = 9'h166 == r_count_34_io_out ? io_r_358_b : _GEN_14137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14139 = 9'h167 == r_count_34_io_out ? io_r_359_b : _GEN_14138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14140 = 9'h168 == r_count_34_io_out ? io_r_360_b : _GEN_14139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14141 = 9'h169 == r_count_34_io_out ? io_r_361_b : _GEN_14140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14142 = 9'h16a == r_count_34_io_out ? io_r_362_b : _GEN_14141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14143 = 9'h16b == r_count_34_io_out ? io_r_363_b : _GEN_14142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14144 = 9'h16c == r_count_34_io_out ? io_r_364_b : _GEN_14143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14145 = 9'h16d == r_count_34_io_out ? io_r_365_b : _GEN_14144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14146 = 9'h16e == r_count_34_io_out ? io_r_366_b : _GEN_14145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14147 = 9'h16f == r_count_34_io_out ? io_r_367_b : _GEN_14146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14148 = 9'h170 == r_count_34_io_out ? io_r_368_b : _GEN_14147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14149 = 9'h171 == r_count_34_io_out ? io_r_369_b : _GEN_14148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14150 = 9'h172 == r_count_34_io_out ? io_r_370_b : _GEN_14149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14151 = 9'h173 == r_count_34_io_out ? io_r_371_b : _GEN_14150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14152 = 9'h174 == r_count_34_io_out ? io_r_372_b : _GEN_14151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14153 = 9'h175 == r_count_34_io_out ? io_r_373_b : _GEN_14152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14154 = 9'h176 == r_count_34_io_out ? io_r_374_b : _GEN_14153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14155 = 9'h177 == r_count_34_io_out ? io_r_375_b : _GEN_14154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14156 = 9'h178 == r_count_34_io_out ? io_r_376_b : _GEN_14155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14157 = 9'h179 == r_count_34_io_out ? io_r_377_b : _GEN_14156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14158 = 9'h17a == r_count_34_io_out ? io_r_378_b : _GEN_14157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14159 = 9'h17b == r_count_34_io_out ? io_r_379_b : _GEN_14158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14160 = 9'h17c == r_count_34_io_out ? io_r_380_b : _GEN_14159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14161 = 9'h17d == r_count_34_io_out ? io_r_381_b : _GEN_14160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14162 = 9'h17e == r_count_34_io_out ? io_r_382_b : _GEN_14161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14163 = 9'h17f == r_count_34_io_out ? io_r_383_b : _GEN_14162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14164 = 9'h180 == r_count_34_io_out ? io_r_384_b : _GEN_14163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14165 = 9'h181 == r_count_34_io_out ? io_r_385_b : _GEN_14164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14166 = 9'h182 == r_count_34_io_out ? io_r_386_b : _GEN_14165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14167 = 9'h183 == r_count_34_io_out ? io_r_387_b : _GEN_14166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14168 = 9'h184 == r_count_34_io_out ? io_r_388_b : _GEN_14167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14169 = 9'h185 == r_count_34_io_out ? io_r_389_b : _GEN_14168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14170 = 9'h186 == r_count_34_io_out ? io_r_390_b : _GEN_14169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14171 = 9'h187 == r_count_34_io_out ? io_r_391_b : _GEN_14170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14172 = 9'h188 == r_count_34_io_out ? io_r_392_b : _GEN_14171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14173 = 9'h189 == r_count_34_io_out ? io_r_393_b : _GEN_14172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14174 = 9'h18a == r_count_34_io_out ? io_r_394_b : _GEN_14173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14175 = 9'h18b == r_count_34_io_out ? io_r_395_b : _GEN_14174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14176 = 9'h18c == r_count_34_io_out ? io_r_396_b : _GEN_14175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14177 = 9'h18d == r_count_34_io_out ? io_r_397_b : _GEN_14176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14178 = 9'h18e == r_count_34_io_out ? io_r_398_b : _GEN_14177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14181 = 9'h1 == r_count_35_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14182 = 9'h2 == r_count_35_io_out ? io_r_2_b : _GEN_14181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14183 = 9'h3 == r_count_35_io_out ? io_r_3_b : _GEN_14182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14184 = 9'h4 == r_count_35_io_out ? io_r_4_b : _GEN_14183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14185 = 9'h5 == r_count_35_io_out ? io_r_5_b : _GEN_14184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14186 = 9'h6 == r_count_35_io_out ? io_r_6_b : _GEN_14185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14187 = 9'h7 == r_count_35_io_out ? io_r_7_b : _GEN_14186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14188 = 9'h8 == r_count_35_io_out ? io_r_8_b : _GEN_14187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14189 = 9'h9 == r_count_35_io_out ? io_r_9_b : _GEN_14188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14190 = 9'ha == r_count_35_io_out ? io_r_10_b : _GEN_14189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14191 = 9'hb == r_count_35_io_out ? io_r_11_b : _GEN_14190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14192 = 9'hc == r_count_35_io_out ? io_r_12_b : _GEN_14191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14193 = 9'hd == r_count_35_io_out ? io_r_13_b : _GEN_14192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14194 = 9'he == r_count_35_io_out ? io_r_14_b : _GEN_14193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14195 = 9'hf == r_count_35_io_out ? io_r_15_b : _GEN_14194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14196 = 9'h10 == r_count_35_io_out ? io_r_16_b : _GEN_14195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14197 = 9'h11 == r_count_35_io_out ? io_r_17_b : _GEN_14196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14198 = 9'h12 == r_count_35_io_out ? io_r_18_b : _GEN_14197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14199 = 9'h13 == r_count_35_io_out ? io_r_19_b : _GEN_14198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14200 = 9'h14 == r_count_35_io_out ? io_r_20_b : _GEN_14199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14201 = 9'h15 == r_count_35_io_out ? io_r_21_b : _GEN_14200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14202 = 9'h16 == r_count_35_io_out ? io_r_22_b : _GEN_14201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14203 = 9'h17 == r_count_35_io_out ? io_r_23_b : _GEN_14202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14204 = 9'h18 == r_count_35_io_out ? io_r_24_b : _GEN_14203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14205 = 9'h19 == r_count_35_io_out ? io_r_25_b : _GEN_14204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14206 = 9'h1a == r_count_35_io_out ? io_r_26_b : _GEN_14205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14207 = 9'h1b == r_count_35_io_out ? io_r_27_b : _GEN_14206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14208 = 9'h1c == r_count_35_io_out ? io_r_28_b : _GEN_14207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14209 = 9'h1d == r_count_35_io_out ? io_r_29_b : _GEN_14208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14210 = 9'h1e == r_count_35_io_out ? io_r_30_b : _GEN_14209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14211 = 9'h1f == r_count_35_io_out ? io_r_31_b : _GEN_14210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14212 = 9'h20 == r_count_35_io_out ? io_r_32_b : _GEN_14211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14213 = 9'h21 == r_count_35_io_out ? io_r_33_b : _GEN_14212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14214 = 9'h22 == r_count_35_io_out ? io_r_34_b : _GEN_14213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14215 = 9'h23 == r_count_35_io_out ? io_r_35_b : _GEN_14214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14216 = 9'h24 == r_count_35_io_out ? io_r_36_b : _GEN_14215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14217 = 9'h25 == r_count_35_io_out ? io_r_37_b : _GEN_14216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14218 = 9'h26 == r_count_35_io_out ? io_r_38_b : _GEN_14217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14219 = 9'h27 == r_count_35_io_out ? io_r_39_b : _GEN_14218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14220 = 9'h28 == r_count_35_io_out ? io_r_40_b : _GEN_14219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14221 = 9'h29 == r_count_35_io_out ? io_r_41_b : _GEN_14220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14222 = 9'h2a == r_count_35_io_out ? io_r_42_b : _GEN_14221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14223 = 9'h2b == r_count_35_io_out ? io_r_43_b : _GEN_14222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14224 = 9'h2c == r_count_35_io_out ? io_r_44_b : _GEN_14223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14225 = 9'h2d == r_count_35_io_out ? io_r_45_b : _GEN_14224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14226 = 9'h2e == r_count_35_io_out ? io_r_46_b : _GEN_14225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14227 = 9'h2f == r_count_35_io_out ? io_r_47_b : _GEN_14226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14228 = 9'h30 == r_count_35_io_out ? io_r_48_b : _GEN_14227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14229 = 9'h31 == r_count_35_io_out ? io_r_49_b : _GEN_14228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14230 = 9'h32 == r_count_35_io_out ? io_r_50_b : _GEN_14229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14231 = 9'h33 == r_count_35_io_out ? io_r_51_b : _GEN_14230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14232 = 9'h34 == r_count_35_io_out ? io_r_52_b : _GEN_14231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14233 = 9'h35 == r_count_35_io_out ? io_r_53_b : _GEN_14232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14234 = 9'h36 == r_count_35_io_out ? io_r_54_b : _GEN_14233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14235 = 9'h37 == r_count_35_io_out ? io_r_55_b : _GEN_14234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14236 = 9'h38 == r_count_35_io_out ? io_r_56_b : _GEN_14235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14237 = 9'h39 == r_count_35_io_out ? io_r_57_b : _GEN_14236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14238 = 9'h3a == r_count_35_io_out ? io_r_58_b : _GEN_14237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14239 = 9'h3b == r_count_35_io_out ? io_r_59_b : _GEN_14238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14240 = 9'h3c == r_count_35_io_out ? io_r_60_b : _GEN_14239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14241 = 9'h3d == r_count_35_io_out ? io_r_61_b : _GEN_14240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14242 = 9'h3e == r_count_35_io_out ? io_r_62_b : _GEN_14241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14243 = 9'h3f == r_count_35_io_out ? io_r_63_b : _GEN_14242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14244 = 9'h40 == r_count_35_io_out ? io_r_64_b : _GEN_14243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14245 = 9'h41 == r_count_35_io_out ? io_r_65_b : _GEN_14244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14246 = 9'h42 == r_count_35_io_out ? io_r_66_b : _GEN_14245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14247 = 9'h43 == r_count_35_io_out ? io_r_67_b : _GEN_14246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14248 = 9'h44 == r_count_35_io_out ? io_r_68_b : _GEN_14247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14249 = 9'h45 == r_count_35_io_out ? io_r_69_b : _GEN_14248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14250 = 9'h46 == r_count_35_io_out ? io_r_70_b : _GEN_14249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14251 = 9'h47 == r_count_35_io_out ? io_r_71_b : _GEN_14250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14252 = 9'h48 == r_count_35_io_out ? io_r_72_b : _GEN_14251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14253 = 9'h49 == r_count_35_io_out ? io_r_73_b : _GEN_14252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14254 = 9'h4a == r_count_35_io_out ? io_r_74_b : _GEN_14253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14255 = 9'h4b == r_count_35_io_out ? io_r_75_b : _GEN_14254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14256 = 9'h4c == r_count_35_io_out ? io_r_76_b : _GEN_14255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14257 = 9'h4d == r_count_35_io_out ? io_r_77_b : _GEN_14256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14258 = 9'h4e == r_count_35_io_out ? io_r_78_b : _GEN_14257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14259 = 9'h4f == r_count_35_io_out ? io_r_79_b : _GEN_14258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14260 = 9'h50 == r_count_35_io_out ? io_r_80_b : _GEN_14259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14261 = 9'h51 == r_count_35_io_out ? io_r_81_b : _GEN_14260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14262 = 9'h52 == r_count_35_io_out ? io_r_82_b : _GEN_14261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14263 = 9'h53 == r_count_35_io_out ? io_r_83_b : _GEN_14262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14264 = 9'h54 == r_count_35_io_out ? io_r_84_b : _GEN_14263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14265 = 9'h55 == r_count_35_io_out ? io_r_85_b : _GEN_14264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14266 = 9'h56 == r_count_35_io_out ? io_r_86_b : _GEN_14265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14267 = 9'h57 == r_count_35_io_out ? io_r_87_b : _GEN_14266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14268 = 9'h58 == r_count_35_io_out ? io_r_88_b : _GEN_14267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14269 = 9'h59 == r_count_35_io_out ? io_r_89_b : _GEN_14268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14270 = 9'h5a == r_count_35_io_out ? io_r_90_b : _GEN_14269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14271 = 9'h5b == r_count_35_io_out ? io_r_91_b : _GEN_14270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14272 = 9'h5c == r_count_35_io_out ? io_r_92_b : _GEN_14271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14273 = 9'h5d == r_count_35_io_out ? io_r_93_b : _GEN_14272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14274 = 9'h5e == r_count_35_io_out ? io_r_94_b : _GEN_14273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14275 = 9'h5f == r_count_35_io_out ? io_r_95_b : _GEN_14274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14276 = 9'h60 == r_count_35_io_out ? io_r_96_b : _GEN_14275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14277 = 9'h61 == r_count_35_io_out ? io_r_97_b : _GEN_14276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14278 = 9'h62 == r_count_35_io_out ? io_r_98_b : _GEN_14277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14279 = 9'h63 == r_count_35_io_out ? io_r_99_b : _GEN_14278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14280 = 9'h64 == r_count_35_io_out ? io_r_100_b : _GEN_14279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14281 = 9'h65 == r_count_35_io_out ? io_r_101_b : _GEN_14280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14282 = 9'h66 == r_count_35_io_out ? io_r_102_b : _GEN_14281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14283 = 9'h67 == r_count_35_io_out ? io_r_103_b : _GEN_14282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14284 = 9'h68 == r_count_35_io_out ? io_r_104_b : _GEN_14283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14285 = 9'h69 == r_count_35_io_out ? io_r_105_b : _GEN_14284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14286 = 9'h6a == r_count_35_io_out ? io_r_106_b : _GEN_14285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14287 = 9'h6b == r_count_35_io_out ? io_r_107_b : _GEN_14286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14288 = 9'h6c == r_count_35_io_out ? io_r_108_b : _GEN_14287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14289 = 9'h6d == r_count_35_io_out ? io_r_109_b : _GEN_14288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14290 = 9'h6e == r_count_35_io_out ? io_r_110_b : _GEN_14289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14291 = 9'h6f == r_count_35_io_out ? io_r_111_b : _GEN_14290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14292 = 9'h70 == r_count_35_io_out ? io_r_112_b : _GEN_14291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14293 = 9'h71 == r_count_35_io_out ? io_r_113_b : _GEN_14292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14294 = 9'h72 == r_count_35_io_out ? io_r_114_b : _GEN_14293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14295 = 9'h73 == r_count_35_io_out ? io_r_115_b : _GEN_14294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14296 = 9'h74 == r_count_35_io_out ? io_r_116_b : _GEN_14295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14297 = 9'h75 == r_count_35_io_out ? io_r_117_b : _GEN_14296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14298 = 9'h76 == r_count_35_io_out ? io_r_118_b : _GEN_14297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14299 = 9'h77 == r_count_35_io_out ? io_r_119_b : _GEN_14298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14300 = 9'h78 == r_count_35_io_out ? io_r_120_b : _GEN_14299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14301 = 9'h79 == r_count_35_io_out ? io_r_121_b : _GEN_14300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14302 = 9'h7a == r_count_35_io_out ? io_r_122_b : _GEN_14301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14303 = 9'h7b == r_count_35_io_out ? io_r_123_b : _GEN_14302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14304 = 9'h7c == r_count_35_io_out ? io_r_124_b : _GEN_14303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14305 = 9'h7d == r_count_35_io_out ? io_r_125_b : _GEN_14304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14306 = 9'h7e == r_count_35_io_out ? io_r_126_b : _GEN_14305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14307 = 9'h7f == r_count_35_io_out ? io_r_127_b : _GEN_14306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14308 = 9'h80 == r_count_35_io_out ? io_r_128_b : _GEN_14307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14309 = 9'h81 == r_count_35_io_out ? io_r_129_b : _GEN_14308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14310 = 9'h82 == r_count_35_io_out ? io_r_130_b : _GEN_14309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14311 = 9'h83 == r_count_35_io_out ? io_r_131_b : _GEN_14310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14312 = 9'h84 == r_count_35_io_out ? io_r_132_b : _GEN_14311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14313 = 9'h85 == r_count_35_io_out ? io_r_133_b : _GEN_14312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14314 = 9'h86 == r_count_35_io_out ? io_r_134_b : _GEN_14313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14315 = 9'h87 == r_count_35_io_out ? io_r_135_b : _GEN_14314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14316 = 9'h88 == r_count_35_io_out ? io_r_136_b : _GEN_14315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14317 = 9'h89 == r_count_35_io_out ? io_r_137_b : _GEN_14316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14318 = 9'h8a == r_count_35_io_out ? io_r_138_b : _GEN_14317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14319 = 9'h8b == r_count_35_io_out ? io_r_139_b : _GEN_14318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14320 = 9'h8c == r_count_35_io_out ? io_r_140_b : _GEN_14319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14321 = 9'h8d == r_count_35_io_out ? io_r_141_b : _GEN_14320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14322 = 9'h8e == r_count_35_io_out ? io_r_142_b : _GEN_14321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14323 = 9'h8f == r_count_35_io_out ? io_r_143_b : _GEN_14322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14324 = 9'h90 == r_count_35_io_out ? io_r_144_b : _GEN_14323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14325 = 9'h91 == r_count_35_io_out ? io_r_145_b : _GEN_14324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14326 = 9'h92 == r_count_35_io_out ? io_r_146_b : _GEN_14325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14327 = 9'h93 == r_count_35_io_out ? io_r_147_b : _GEN_14326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14328 = 9'h94 == r_count_35_io_out ? io_r_148_b : _GEN_14327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14329 = 9'h95 == r_count_35_io_out ? io_r_149_b : _GEN_14328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14330 = 9'h96 == r_count_35_io_out ? io_r_150_b : _GEN_14329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14331 = 9'h97 == r_count_35_io_out ? io_r_151_b : _GEN_14330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14332 = 9'h98 == r_count_35_io_out ? io_r_152_b : _GEN_14331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14333 = 9'h99 == r_count_35_io_out ? io_r_153_b : _GEN_14332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14334 = 9'h9a == r_count_35_io_out ? io_r_154_b : _GEN_14333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14335 = 9'h9b == r_count_35_io_out ? io_r_155_b : _GEN_14334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14336 = 9'h9c == r_count_35_io_out ? io_r_156_b : _GEN_14335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14337 = 9'h9d == r_count_35_io_out ? io_r_157_b : _GEN_14336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14338 = 9'h9e == r_count_35_io_out ? io_r_158_b : _GEN_14337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14339 = 9'h9f == r_count_35_io_out ? io_r_159_b : _GEN_14338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14340 = 9'ha0 == r_count_35_io_out ? io_r_160_b : _GEN_14339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14341 = 9'ha1 == r_count_35_io_out ? io_r_161_b : _GEN_14340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14342 = 9'ha2 == r_count_35_io_out ? io_r_162_b : _GEN_14341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14343 = 9'ha3 == r_count_35_io_out ? io_r_163_b : _GEN_14342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14344 = 9'ha4 == r_count_35_io_out ? io_r_164_b : _GEN_14343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14345 = 9'ha5 == r_count_35_io_out ? io_r_165_b : _GEN_14344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14346 = 9'ha6 == r_count_35_io_out ? io_r_166_b : _GEN_14345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14347 = 9'ha7 == r_count_35_io_out ? io_r_167_b : _GEN_14346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14348 = 9'ha8 == r_count_35_io_out ? io_r_168_b : _GEN_14347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14349 = 9'ha9 == r_count_35_io_out ? io_r_169_b : _GEN_14348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14350 = 9'haa == r_count_35_io_out ? io_r_170_b : _GEN_14349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14351 = 9'hab == r_count_35_io_out ? io_r_171_b : _GEN_14350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14352 = 9'hac == r_count_35_io_out ? io_r_172_b : _GEN_14351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14353 = 9'had == r_count_35_io_out ? io_r_173_b : _GEN_14352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14354 = 9'hae == r_count_35_io_out ? io_r_174_b : _GEN_14353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14355 = 9'haf == r_count_35_io_out ? io_r_175_b : _GEN_14354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14356 = 9'hb0 == r_count_35_io_out ? io_r_176_b : _GEN_14355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14357 = 9'hb1 == r_count_35_io_out ? io_r_177_b : _GEN_14356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14358 = 9'hb2 == r_count_35_io_out ? io_r_178_b : _GEN_14357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14359 = 9'hb3 == r_count_35_io_out ? io_r_179_b : _GEN_14358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14360 = 9'hb4 == r_count_35_io_out ? io_r_180_b : _GEN_14359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14361 = 9'hb5 == r_count_35_io_out ? io_r_181_b : _GEN_14360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14362 = 9'hb6 == r_count_35_io_out ? io_r_182_b : _GEN_14361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14363 = 9'hb7 == r_count_35_io_out ? io_r_183_b : _GEN_14362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14364 = 9'hb8 == r_count_35_io_out ? io_r_184_b : _GEN_14363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14365 = 9'hb9 == r_count_35_io_out ? io_r_185_b : _GEN_14364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14366 = 9'hba == r_count_35_io_out ? io_r_186_b : _GEN_14365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14367 = 9'hbb == r_count_35_io_out ? io_r_187_b : _GEN_14366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14368 = 9'hbc == r_count_35_io_out ? io_r_188_b : _GEN_14367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14369 = 9'hbd == r_count_35_io_out ? io_r_189_b : _GEN_14368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14370 = 9'hbe == r_count_35_io_out ? io_r_190_b : _GEN_14369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14371 = 9'hbf == r_count_35_io_out ? io_r_191_b : _GEN_14370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14372 = 9'hc0 == r_count_35_io_out ? io_r_192_b : _GEN_14371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14373 = 9'hc1 == r_count_35_io_out ? io_r_193_b : _GEN_14372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14374 = 9'hc2 == r_count_35_io_out ? io_r_194_b : _GEN_14373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14375 = 9'hc3 == r_count_35_io_out ? io_r_195_b : _GEN_14374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14376 = 9'hc4 == r_count_35_io_out ? io_r_196_b : _GEN_14375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14377 = 9'hc5 == r_count_35_io_out ? io_r_197_b : _GEN_14376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14378 = 9'hc6 == r_count_35_io_out ? io_r_198_b : _GEN_14377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14379 = 9'hc7 == r_count_35_io_out ? io_r_199_b : _GEN_14378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14380 = 9'hc8 == r_count_35_io_out ? io_r_200_b : _GEN_14379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14381 = 9'hc9 == r_count_35_io_out ? io_r_201_b : _GEN_14380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14382 = 9'hca == r_count_35_io_out ? io_r_202_b : _GEN_14381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14383 = 9'hcb == r_count_35_io_out ? io_r_203_b : _GEN_14382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14384 = 9'hcc == r_count_35_io_out ? io_r_204_b : _GEN_14383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14385 = 9'hcd == r_count_35_io_out ? io_r_205_b : _GEN_14384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14386 = 9'hce == r_count_35_io_out ? io_r_206_b : _GEN_14385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14387 = 9'hcf == r_count_35_io_out ? io_r_207_b : _GEN_14386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14388 = 9'hd0 == r_count_35_io_out ? io_r_208_b : _GEN_14387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14389 = 9'hd1 == r_count_35_io_out ? io_r_209_b : _GEN_14388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14390 = 9'hd2 == r_count_35_io_out ? io_r_210_b : _GEN_14389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14391 = 9'hd3 == r_count_35_io_out ? io_r_211_b : _GEN_14390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14392 = 9'hd4 == r_count_35_io_out ? io_r_212_b : _GEN_14391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14393 = 9'hd5 == r_count_35_io_out ? io_r_213_b : _GEN_14392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14394 = 9'hd6 == r_count_35_io_out ? io_r_214_b : _GEN_14393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14395 = 9'hd7 == r_count_35_io_out ? io_r_215_b : _GEN_14394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14396 = 9'hd8 == r_count_35_io_out ? io_r_216_b : _GEN_14395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14397 = 9'hd9 == r_count_35_io_out ? io_r_217_b : _GEN_14396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14398 = 9'hda == r_count_35_io_out ? io_r_218_b : _GEN_14397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14399 = 9'hdb == r_count_35_io_out ? io_r_219_b : _GEN_14398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14400 = 9'hdc == r_count_35_io_out ? io_r_220_b : _GEN_14399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14401 = 9'hdd == r_count_35_io_out ? io_r_221_b : _GEN_14400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14402 = 9'hde == r_count_35_io_out ? io_r_222_b : _GEN_14401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14403 = 9'hdf == r_count_35_io_out ? io_r_223_b : _GEN_14402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14404 = 9'he0 == r_count_35_io_out ? io_r_224_b : _GEN_14403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14405 = 9'he1 == r_count_35_io_out ? io_r_225_b : _GEN_14404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14406 = 9'he2 == r_count_35_io_out ? io_r_226_b : _GEN_14405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14407 = 9'he3 == r_count_35_io_out ? io_r_227_b : _GEN_14406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14408 = 9'he4 == r_count_35_io_out ? io_r_228_b : _GEN_14407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14409 = 9'he5 == r_count_35_io_out ? io_r_229_b : _GEN_14408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14410 = 9'he6 == r_count_35_io_out ? io_r_230_b : _GEN_14409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14411 = 9'he7 == r_count_35_io_out ? io_r_231_b : _GEN_14410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14412 = 9'he8 == r_count_35_io_out ? io_r_232_b : _GEN_14411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14413 = 9'he9 == r_count_35_io_out ? io_r_233_b : _GEN_14412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14414 = 9'hea == r_count_35_io_out ? io_r_234_b : _GEN_14413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14415 = 9'heb == r_count_35_io_out ? io_r_235_b : _GEN_14414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14416 = 9'hec == r_count_35_io_out ? io_r_236_b : _GEN_14415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14417 = 9'hed == r_count_35_io_out ? io_r_237_b : _GEN_14416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14418 = 9'hee == r_count_35_io_out ? io_r_238_b : _GEN_14417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14419 = 9'hef == r_count_35_io_out ? io_r_239_b : _GEN_14418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14420 = 9'hf0 == r_count_35_io_out ? io_r_240_b : _GEN_14419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14421 = 9'hf1 == r_count_35_io_out ? io_r_241_b : _GEN_14420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14422 = 9'hf2 == r_count_35_io_out ? io_r_242_b : _GEN_14421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14423 = 9'hf3 == r_count_35_io_out ? io_r_243_b : _GEN_14422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14424 = 9'hf4 == r_count_35_io_out ? io_r_244_b : _GEN_14423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14425 = 9'hf5 == r_count_35_io_out ? io_r_245_b : _GEN_14424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14426 = 9'hf6 == r_count_35_io_out ? io_r_246_b : _GEN_14425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14427 = 9'hf7 == r_count_35_io_out ? io_r_247_b : _GEN_14426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14428 = 9'hf8 == r_count_35_io_out ? io_r_248_b : _GEN_14427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14429 = 9'hf9 == r_count_35_io_out ? io_r_249_b : _GEN_14428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14430 = 9'hfa == r_count_35_io_out ? io_r_250_b : _GEN_14429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14431 = 9'hfb == r_count_35_io_out ? io_r_251_b : _GEN_14430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14432 = 9'hfc == r_count_35_io_out ? io_r_252_b : _GEN_14431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14433 = 9'hfd == r_count_35_io_out ? io_r_253_b : _GEN_14432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14434 = 9'hfe == r_count_35_io_out ? io_r_254_b : _GEN_14433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14435 = 9'hff == r_count_35_io_out ? io_r_255_b : _GEN_14434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14436 = 9'h100 == r_count_35_io_out ? io_r_256_b : _GEN_14435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14437 = 9'h101 == r_count_35_io_out ? io_r_257_b : _GEN_14436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14438 = 9'h102 == r_count_35_io_out ? io_r_258_b : _GEN_14437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14439 = 9'h103 == r_count_35_io_out ? io_r_259_b : _GEN_14438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14440 = 9'h104 == r_count_35_io_out ? io_r_260_b : _GEN_14439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14441 = 9'h105 == r_count_35_io_out ? io_r_261_b : _GEN_14440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14442 = 9'h106 == r_count_35_io_out ? io_r_262_b : _GEN_14441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14443 = 9'h107 == r_count_35_io_out ? io_r_263_b : _GEN_14442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14444 = 9'h108 == r_count_35_io_out ? io_r_264_b : _GEN_14443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14445 = 9'h109 == r_count_35_io_out ? io_r_265_b : _GEN_14444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14446 = 9'h10a == r_count_35_io_out ? io_r_266_b : _GEN_14445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14447 = 9'h10b == r_count_35_io_out ? io_r_267_b : _GEN_14446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14448 = 9'h10c == r_count_35_io_out ? io_r_268_b : _GEN_14447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14449 = 9'h10d == r_count_35_io_out ? io_r_269_b : _GEN_14448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14450 = 9'h10e == r_count_35_io_out ? io_r_270_b : _GEN_14449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14451 = 9'h10f == r_count_35_io_out ? io_r_271_b : _GEN_14450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14452 = 9'h110 == r_count_35_io_out ? io_r_272_b : _GEN_14451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14453 = 9'h111 == r_count_35_io_out ? io_r_273_b : _GEN_14452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14454 = 9'h112 == r_count_35_io_out ? io_r_274_b : _GEN_14453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14455 = 9'h113 == r_count_35_io_out ? io_r_275_b : _GEN_14454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14456 = 9'h114 == r_count_35_io_out ? io_r_276_b : _GEN_14455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14457 = 9'h115 == r_count_35_io_out ? io_r_277_b : _GEN_14456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14458 = 9'h116 == r_count_35_io_out ? io_r_278_b : _GEN_14457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14459 = 9'h117 == r_count_35_io_out ? io_r_279_b : _GEN_14458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14460 = 9'h118 == r_count_35_io_out ? io_r_280_b : _GEN_14459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14461 = 9'h119 == r_count_35_io_out ? io_r_281_b : _GEN_14460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14462 = 9'h11a == r_count_35_io_out ? io_r_282_b : _GEN_14461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14463 = 9'h11b == r_count_35_io_out ? io_r_283_b : _GEN_14462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14464 = 9'h11c == r_count_35_io_out ? io_r_284_b : _GEN_14463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14465 = 9'h11d == r_count_35_io_out ? io_r_285_b : _GEN_14464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14466 = 9'h11e == r_count_35_io_out ? io_r_286_b : _GEN_14465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14467 = 9'h11f == r_count_35_io_out ? io_r_287_b : _GEN_14466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14468 = 9'h120 == r_count_35_io_out ? io_r_288_b : _GEN_14467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14469 = 9'h121 == r_count_35_io_out ? io_r_289_b : _GEN_14468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14470 = 9'h122 == r_count_35_io_out ? io_r_290_b : _GEN_14469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14471 = 9'h123 == r_count_35_io_out ? io_r_291_b : _GEN_14470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14472 = 9'h124 == r_count_35_io_out ? io_r_292_b : _GEN_14471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14473 = 9'h125 == r_count_35_io_out ? io_r_293_b : _GEN_14472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14474 = 9'h126 == r_count_35_io_out ? io_r_294_b : _GEN_14473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14475 = 9'h127 == r_count_35_io_out ? io_r_295_b : _GEN_14474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14476 = 9'h128 == r_count_35_io_out ? io_r_296_b : _GEN_14475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14477 = 9'h129 == r_count_35_io_out ? io_r_297_b : _GEN_14476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14478 = 9'h12a == r_count_35_io_out ? io_r_298_b : _GEN_14477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14479 = 9'h12b == r_count_35_io_out ? io_r_299_b : _GEN_14478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14480 = 9'h12c == r_count_35_io_out ? io_r_300_b : _GEN_14479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14481 = 9'h12d == r_count_35_io_out ? io_r_301_b : _GEN_14480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14482 = 9'h12e == r_count_35_io_out ? io_r_302_b : _GEN_14481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14483 = 9'h12f == r_count_35_io_out ? io_r_303_b : _GEN_14482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14484 = 9'h130 == r_count_35_io_out ? io_r_304_b : _GEN_14483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14485 = 9'h131 == r_count_35_io_out ? io_r_305_b : _GEN_14484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14486 = 9'h132 == r_count_35_io_out ? io_r_306_b : _GEN_14485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14487 = 9'h133 == r_count_35_io_out ? io_r_307_b : _GEN_14486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14488 = 9'h134 == r_count_35_io_out ? io_r_308_b : _GEN_14487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14489 = 9'h135 == r_count_35_io_out ? io_r_309_b : _GEN_14488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14490 = 9'h136 == r_count_35_io_out ? io_r_310_b : _GEN_14489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14491 = 9'h137 == r_count_35_io_out ? io_r_311_b : _GEN_14490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14492 = 9'h138 == r_count_35_io_out ? io_r_312_b : _GEN_14491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14493 = 9'h139 == r_count_35_io_out ? io_r_313_b : _GEN_14492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14494 = 9'h13a == r_count_35_io_out ? io_r_314_b : _GEN_14493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14495 = 9'h13b == r_count_35_io_out ? io_r_315_b : _GEN_14494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14496 = 9'h13c == r_count_35_io_out ? io_r_316_b : _GEN_14495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14497 = 9'h13d == r_count_35_io_out ? io_r_317_b : _GEN_14496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14498 = 9'h13e == r_count_35_io_out ? io_r_318_b : _GEN_14497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14499 = 9'h13f == r_count_35_io_out ? io_r_319_b : _GEN_14498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14500 = 9'h140 == r_count_35_io_out ? io_r_320_b : _GEN_14499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14501 = 9'h141 == r_count_35_io_out ? io_r_321_b : _GEN_14500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14502 = 9'h142 == r_count_35_io_out ? io_r_322_b : _GEN_14501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14503 = 9'h143 == r_count_35_io_out ? io_r_323_b : _GEN_14502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14504 = 9'h144 == r_count_35_io_out ? io_r_324_b : _GEN_14503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14505 = 9'h145 == r_count_35_io_out ? io_r_325_b : _GEN_14504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14506 = 9'h146 == r_count_35_io_out ? io_r_326_b : _GEN_14505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14507 = 9'h147 == r_count_35_io_out ? io_r_327_b : _GEN_14506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14508 = 9'h148 == r_count_35_io_out ? io_r_328_b : _GEN_14507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14509 = 9'h149 == r_count_35_io_out ? io_r_329_b : _GEN_14508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14510 = 9'h14a == r_count_35_io_out ? io_r_330_b : _GEN_14509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14511 = 9'h14b == r_count_35_io_out ? io_r_331_b : _GEN_14510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14512 = 9'h14c == r_count_35_io_out ? io_r_332_b : _GEN_14511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14513 = 9'h14d == r_count_35_io_out ? io_r_333_b : _GEN_14512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14514 = 9'h14e == r_count_35_io_out ? io_r_334_b : _GEN_14513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14515 = 9'h14f == r_count_35_io_out ? io_r_335_b : _GEN_14514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14516 = 9'h150 == r_count_35_io_out ? io_r_336_b : _GEN_14515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14517 = 9'h151 == r_count_35_io_out ? io_r_337_b : _GEN_14516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14518 = 9'h152 == r_count_35_io_out ? io_r_338_b : _GEN_14517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14519 = 9'h153 == r_count_35_io_out ? io_r_339_b : _GEN_14518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14520 = 9'h154 == r_count_35_io_out ? io_r_340_b : _GEN_14519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14521 = 9'h155 == r_count_35_io_out ? io_r_341_b : _GEN_14520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14522 = 9'h156 == r_count_35_io_out ? io_r_342_b : _GEN_14521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14523 = 9'h157 == r_count_35_io_out ? io_r_343_b : _GEN_14522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14524 = 9'h158 == r_count_35_io_out ? io_r_344_b : _GEN_14523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14525 = 9'h159 == r_count_35_io_out ? io_r_345_b : _GEN_14524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14526 = 9'h15a == r_count_35_io_out ? io_r_346_b : _GEN_14525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14527 = 9'h15b == r_count_35_io_out ? io_r_347_b : _GEN_14526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14528 = 9'h15c == r_count_35_io_out ? io_r_348_b : _GEN_14527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14529 = 9'h15d == r_count_35_io_out ? io_r_349_b : _GEN_14528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14530 = 9'h15e == r_count_35_io_out ? io_r_350_b : _GEN_14529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14531 = 9'h15f == r_count_35_io_out ? io_r_351_b : _GEN_14530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14532 = 9'h160 == r_count_35_io_out ? io_r_352_b : _GEN_14531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14533 = 9'h161 == r_count_35_io_out ? io_r_353_b : _GEN_14532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14534 = 9'h162 == r_count_35_io_out ? io_r_354_b : _GEN_14533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14535 = 9'h163 == r_count_35_io_out ? io_r_355_b : _GEN_14534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14536 = 9'h164 == r_count_35_io_out ? io_r_356_b : _GEN_14535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14537 = 9'h165 == r_count_35_io_out ? io_r_357_b : _GEN_14536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14538 = 9'h166 == r_count_35_io_out ? io_r_358_b : _GEN_14537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14539 = 9'h167 == r_count_35_io_out ? io_r_359_b : _GEN_14538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14540 = 9'h168 == r_count_35_io_out ? io_r_360_b : _GEN_14539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14541 = 9'h169 == r_count_35_io_out ? io_r_361_b : _GEN_14540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14542 = 9'h16a == r_count_35_io_out ? io_r_362_b : _GEN_14541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14543 = 9'h16b == r_count_35_io_out ? io_r_363_b : _GEN_14542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14544 = 9'h16c == r_count_35_io_out ? io_r_364_b : _GEN_14543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14545 = 9'h16d == r_count_35_io_out ? io_r_365_b : _GEN_14544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14546 = 9'h16e == r_count_35_io_out ? io_r_366_b : _GEN_14545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14547 = 9'h16f == r_count_35_io_out ? io_r_367_b : _GEN_14546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14548 = 9'h170 == r_count_35_io_out ? io_r_368_b : _GEN_14547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14549 = 9'h171 == r_count_35_io_out ? io_r_369_b : _GEN_14548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14550 = 9'h172 == r_count_35_io_out ? io_r_370_b : _GEN_14549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14551 = 9'h173 == r_count_35_io_out ? io_r_371_b : _GEN_14550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14552 = 9'h174 == r_count_35_io_out ? io_r_372_b : _GEN_14551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14553 = 9'h175 == r_count_35_io_out ? io_r_373_b : _GEN_14552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14554 = 9'h176 == r_count_35_io_out ? io_r_374_b : _GEN_14553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14555 = 9'h177 == r_count_35_io_out ? io_r_375_b : _GEN_14554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14556 = 9'h178 == r_count_35_io_out ? io_r_376_b : _GEN_14555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14557 = 9'h179 == r_count_35_io_out ? io_r_377_b : _GEN_14556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14558 = 9'h17a == r_count_35_io_out ? io_r_378_b : _GEN_14557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14559 = 9'h17b == r_count_35_io_out ? io_r_379_b : _GEN_14558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14560 = 9'h17c == r_count_35_io_out ? io_r_380_b : _GEN_14559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14561 = 9'h17d == r_count_35_io_out ? io_r_381_b : _GEN_14560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14562 = 9'h17e == r_count_35_io_out ? io_r_382_b : _GEN_14561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14563 = 9'h17f == r_count_35_io_out ? io_r_383_b : _GEN_14562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14564 = 9'h180 == r_count_35_io_out ? io_r_384_b : _GEN_14563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14565 = 9'h181 == r_count_35_io_out ? io_r_385_b : _GEN_14564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14566 = 9'h182 == r_count_35_io_out ? io_r_386_b : _GEN_14565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14567 = 9'h183 == r_count_35_io_out ? io_r_387_b : _GEN_14566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14568 = 9'h184 == r_count_35_io_out ? io_r_388_b : _GEN_14567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14569 = 9'h185 == r_count_35_io_out ? io_r_389_b : _GEN_14568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14570 = 9'h186 == r_count_35_io_out ? io_r_390_b : _GEN_14569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14571 = 9'h187 == r_count_35_io_out ? io_r_391_b : _GEN_14570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14572 = 9'h188 == r_count_35_io_out ? io_r_392_b : _GEN_14571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14573 = 9'h189 == r_count_35_io_out ? io_r_393_b : _GEN_14572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14574 = 9'h18a == r_count_35_io_out ? io_r_394_b : _GEN_14573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14575 = 9'h18b == r_count_35_io_out ? io_r_395_b : _GEN_14574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14576 = 9'h18c == r_count_35_io_out ? io_r_396_b : _GEN_14575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14577 = 9'h18d == r_count_35_io_out ? io_r_397_b : _GEN_14576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14578 = 9'h18e == r_count_35_io_out ? io_r_398_b : _GEN_14577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14581 = 9'h1 == r_count_36_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14582 = 9'h2 == r_count_36_io_out ? io_r_2_b : _GEN_14581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14583 = 9'h3 == r_count_36_io_out ? io_r_3_b : _GEN_14582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14584 = 9'h4 == r_count_36_io_out ? io_r_4_b : _GEN_14583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14585 = 9'h5 == r_count_36_io_out ? io_r_5_b : _GEN_14584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14586 = 9'h6 == r_count_36_io_out ? io_r_6_b : _GEN_14585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14587 = 9'h7 == r_count_36_io_out ? io_r_7_b : _GEN_14586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14588 = 9'h8 == r_count_36_io_out ? io_r_8_b : _GEN_14587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14589 = 9'h9 == r_count_36_io_out ? io_r_9_b : _GEN_14588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14590 = 9'ha == r_count_36_io_out ? io_r_10_b : _GEN_14589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14591 = 9'hb == r_count_36_io_out ? io_r_11_b : _GEN_14590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14592 = 9'hc == r_count_36_io_out ? io_r_12_b : _GEN_14591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14593 = 9'hd == r_count_36_io_out ? io_r_13_b : _GEN_14592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14594 = 9'he == r_count_36_io_out ? io_r_14_b : _GEN_14593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14595 = 9'hf == r_count_36_io_out ? io_r_15_b : _GEN_14594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14596 = 9'h10 == r_count_36_io_out ? io_r_16_b : _GEN_14595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14597 = 9'h11 == r_count_36_io_out ? io_r_17_b : _GEN_14596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14598 = 9'h12 == r_count_36_io_out ? io_r_18_b : _GEN_14597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14599 = 9'h13 == r_count_36_io_out ? io_r_19_b : _GEN_14598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14600 = 9'h14 == r_count_36_io_out ? io_r_20_b : _GEN_14599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14601 = 9'h15 == r_count_36_io_out ? io_r_21_b : _GEN_14600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14602 = 9'h16 == r_count_36_io_out ? io_r_22_b : _GEN_14601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14603 = 9'h17 == r_count_36_io_out ? io_r_23_b : _GEN_14602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14604 = 9'h18 == r_count_36_io_out ? io_r_24_b : _GEN_14603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14605 = 9'h19 == r_count_36_io_out ? io_r_25_b : _GEN_14604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14606 = 9'h1a == r_count_36_io_out ? io_r_26_b : _GEN_14605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14607 = 9'h1b == r_count_36_io_out ? io_r_27_b : _GEN_14606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14608 = 9'h1c == r_count_36_io_out ? io_r_28_b : _GEN_14607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14609 = 9'h1d == r_count_36_io_out ? io_r_29_b : _GEN_14608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14610 = 9'h1e == r_count_36_io_out ? io_r_30_b : _GEN_14609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14611 = 9'h1f == r_count_36_io_out ? io_r_31_b : _GEN_14610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14612 = 9'h20 == r_count_36_io_out ? io_r_32_b : _GEN_14611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14613 = 9'h21 == r_count_36_io_out ? io_r_33_b : _GEN_14612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14614 = 9'h22 == r_count_36_io_out ? io_r_34_b : _GEN_14613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14615 = 9'h23 == r_count_36_io_out ? io_r_35_b : _GEN_14614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14616 = 9'h24 == r_count_36_io_out ? io_r_36_b : _GEN_14615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14617 = 9'h25 == r_count_36_io_out ? io_r_37_b : _GEN_14616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14618 = 9'h26 == r_count_36_io_out ? io_r_38_b : _GEN_14617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14619 = 9'h27 == r_count_36_io_out ? io_r_39_b : _GEN_14618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14620 = 9'h28 == r_count_36_io_out ? io_r_40_b : _GEN_14619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14621 = 9'h29 == r_count_36_io_out ? io_r_41_b : _GEN_14620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14622 = 9'h2a == r_count_36_io_out ? io_r_42_b : _GEN_14621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14623 = 9'h2b == r_count_36_io_out ? io_r_43_b : _GEN_14622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14624 = 9'h2c == r_count_36_io_out ? io_r_44_b : _GEN_14623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14625 = 9'h2d == r_count_36_io_out ? io_r_45_b : _GEN_14624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14626 = 9'h2e == r_count_36_io_out ? io_r_46_b : _GEN_14625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14627 = 9'h2f == r_count_36_io_out ? io_r_47_b : _GEN_14626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14628 = 9'h30 == r_count_36_io_out ? io_r_48_b : _GEN_14627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14629 = 9'h31 == r_count_36_io_out ? io_r_49_b : _GEN_14628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14630 = 9'h32 == r_count_36_io_out ? io_r_50_b : _GEN_14629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14631 = 9'h33 == r_count_36_io_out ? io_r_51_b : _GEN_14630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14632 = 9'h34 == r_count_36_io_out ? io_r_52_b : _GEN_14631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14633 = 9'h35 == r_count_36_io_out ? io_r_53_b : _GEN_14632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14634 = 9'h36 == r_count_36_io_out ? io_r_54_b : _GEN_14633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14635 = 9'h37 == r_count_36_io_out ? io_r_55_b : _GEN_14634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14636 = 9'h38 == r_count_36_io_out ? io_r_56_b : _GEN_14635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14637 = 9'h39 == r_count_36_io_out ? io_r_57_b : _GEN_14636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14638 = 9'h3a == r_count_36_io_out ? io_r_58_b : _GEN_14637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14639 = 9'h3b == r_count_36_io_out ? io_r_59_b : _GEN_14638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14640 = 9'h3c == r_count_36_io_out ? io_r_60_b : _GEN_14639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14641 = 9'h3d == r_count_36_io_out ? io_r_61_b : _GEN_14640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14642 = 9'h3e == r_count_36_io_out ? io_r_62_b : _GEN_14641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14643 = 9'h3f == r_count_36_io_out ? io_r_63_b : _GEN_14642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14644 = 9'h40 == r_count_36_io_out ? io_r_64_b : _GEN_14643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14645 = 9'h41 == r_count_36_io_out ? io_r_65_b : _GEN_14644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14646 = 9'h42 == r_count_36_io_out ? io_r_66_b : _GEN_14645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14647 = 9'h43 == r_count_36_io_out ? io_r_67_b : _GEN_14646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14648 = 9'h44 == r_count_36_io_out ? io_r_68_b : _GEN_14647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14649 = 9'h45 == r_count_36_io_out ? io_r_69_b : _GEN_14648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14650 = 9'h46 == r_count_36_io_out ? io_r_70_b : _GEN_14649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14651 = 9'h47 == r_count_36_io_out ? io_r_71_b : _GEN_14650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14652 = 9'h48 == r_count_36_io_out ? io_r_72_b : _GEN_14651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14653 = 9'h49 == r_count_36_io_out ? io_r_73_b : _GEN_14652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14654 = 9'h4a == r_count_36_io_out ? io_r_74_b : _GEN_14653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14655 = 9'h4b == r_count_36_io_out ? io_r_75_b : _GEN_14654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14656 = 9'h4c == r_count_36_io_out ? io_r_76_b : _GEN_14655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14657 = 9'h4d == r_count_36_io_out ? io_r_77_b : _GEN_14656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14658 = 9'h4e == r_count_36_io_out ? io_r_78_b : _GEN_14657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14659 = 9'h4f == r_count_36_io_out ? io_r_79_b : _GEN_14658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14660 = 9'h50 == r_count_36_io_out ? io_r_80_b : _GEN_14659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14661 = 9'h51 == r_count_36_io_out ? io_r_81_b : _GEN_14660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14662 = 9'h52 == r_count_36_io_out ? io_r_82_b : _GEN_14661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14663 = 9'h53 == r_count_36_io_out ? io_r_83_b : _GEN_14662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14664 = 9'h54 == r_count_36_io_out ? io_r_84_b : _GEN_14663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14665 = 9'h55 == r_count_36_io_out ? io_r_85_b : _GEN_14664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14666 = 9'h56 == r_count_36_io_out ? io_r_86_b : _GEN_14665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14667 = 9'h57 == r_count_36_io_out ? io_r_87_b : _GEN_14666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14668 = 9'h58 == r_count_36_io_out ? io_r_88_b : _GEN_14667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14669 = 9'h59 == r_count_36_io_out ? io_r_89_b : _GEN_14668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14670 = 9'h5a == r_count_36_io_out ? io_r_90_b : _GEN_14669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14671 = 9'h5b == r_count_36_io_out ? io_r_91_b : _GEN_14670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14672 = 9'h5c == r_count_36_io_out ? io_r_92_b : _GEN_14671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14673 = 9'h5d == r_count_36_io_out ? io_r_93_b : _GEN_14672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14674 = 9'h5e == r_count_36_io_out ? io_r_94_b : _GEN_14673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14675 = 9'h5f == r_count_36_io_out ? io_r_95_b : _GEN_14674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14676 = 9'h60 == r_count_36_io_out ? io_r_96_b : _GEN_14675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14677 = 9'h61 == r_count_36_io_out ? io_r_97_b : _GEN_14676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14678 = 9'h62 == r_count_36_io_out ? io_r_98_b : _GEN_14677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14679 = 9'h63 == r_count_36_io_out ? io_r_99_b : _GEN_14678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14680 = 9'h64 == r_count_36_io_out ? io_r_100_b : _GEN_14679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14681 = 9'h65 == r_count_36_io_out ? io_r_101_b : _GEN_14680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14682 = 9'h66 == r_count_36_io_out ? io_r_102_b : _GEN_14681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14683 = 9'h67 == r_count_36_io_out ? io_r_103_b : _GEN_14682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14684 = 9'h68 == r_count_36_io_out ? io_r_104_b : _GEN_14683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14685 = 9'h69 == r_count_36_io_out ? io_r_105_b : _GEN_14684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14686 = 9'h6a == r_count_36_io_out ? io_r_106_b : _GEN_14685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14687 = 9'h6b == r_count_36_io_out ? io_r_107_b : _GEN_14686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14688 = 9'h6c == r_count_36_io_out ? io_r_108_b : _GEN_14687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14689 = 9'h6d == r_count_36_io_out ? io_r_109_b : _GEN_14688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14690 = 9'h6e == r_count_36_io_out ? io_r_110_b : _GEN_14689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14691 = 9'h6f == r_count_36_io_out ? io_r_111_b : _GEN_14690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14692 = 9'h70 == r_count_36_io_out ? io_r_112_b : _GEN_14691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14693 = 9'h71 == r_count_36_io_out ? io_r_113_b : _GEN_14692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14694 = 9'h72 == r_count_36_io_out ? io_r_114_b : _GEN_14693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14695 = 9'h73 == r_count_36_io_out ? io_r_115_b : _GEN_14694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14696 = 9'h74 == r_count_36_io_out ? io_r_116_b : _GEN_14695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14697 = 9'h75 == r_count_36_io_out ? io_r_117_b : _GEN_14696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14698 = 9'h76 == r_count_36_io_out ? io_r_118_b : _GEN_14697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14699 = 9'h77 == r_count_36_io_out ? io_r_119_b : _GEN_14698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14700 = 9'h78 == r_count_36_io_out ? io_r_120_b : _GEN_14699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14701 = 9'h79 == r_count_36_io_out ? io_r_121_b : _GEN_14700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14702 = 9'h7a == r_count_36_io_out ? io_r_122_b : _GEN_14701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14703 = 9'h7b == r_count_36_io_out ? io_r_123_b : _GEN_14702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14704 = 9'h7c == r_count_36_io_out ? io_r_124_b : _GEN_14703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14705 = 9'h7d == r_count_36_io_out ? io_r_125_b : _GEN_14704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14706 = 9'h7e == r_count_36_io_out ? io_r_126_b : _GEN_14705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14707 = 9'h7f == r_count_36_io_out ? io_r_127_b : _GEN_14706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14708 = 9'h80 == r_count_36_io_out ? io_r_128_b : _GEN_14707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14709 = 9'h81 == r_count_36_io_out ? io_r_129_b : _GEN_14708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14710 = 9'h82 == r_count_36_io_out ? io_r_130_b : _GEN_14709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14711 = 9'h83 == r_count_36_io_out ? io_r_131_b : _GEN_14710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14712 = 9'h84 == r_count_36_io_out ? io_r_132_b : _GEN_14711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14713 = 9'h85 == r_count_36_io_out ? io_r_133_b : _GEN_14712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14714 = 9'h86 == r_count_36_io_out ? io_r_134_b : _GEN_14713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14715 = 9'h87 == r_count_36_io_out ? io_r_135_b : _GEN_14714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14716 = 9'h88 == r_count_36_io_out ? io_r_136_b : _GEN_14715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14717 = 9'h89 == r_count_36_io_out ? io_r_137_b : _GEN_14716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14718 = 9'h8a == r_count_36_io_out ? io_r_138_b : _GEN_14717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14719 = 9'h8b == r_count_36_io_out ? io_r_139_b : _GEN_14718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14720 = 9'h8c == r_count_36_io_out ? io_r_140_b : _GEN_14719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14721 = 9'h8d == r_count_36_io_out ? io_r_141_b : _GEN_14720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14722 = 9'h8e == r_count_36_io_out ? io_r_142_b : _GEN_14721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14723 = 9'h8f == r_count_36_io_out ? io_r_143_b : _GEN_14722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14724 = 9'h90 == r_count_36_io_out ? io_r_144_b : _GEN_14723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14725 = 9'h91 == r_count_36_io_out ? io_r_145_b : _GEN_14724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14726 = 9'h92 == r_count_36_io_out ? io_r_146_b : _GEN_14725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14727 = 9'h93 == r_count_36_io_out ? io_r_147_b : _GEN_14726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14728 = 9'h94 == r_count_36_io_out ? io_r_148_b : _GEN_14727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14729 = 9'h95 == r_count_36_io_out ? io_r_149_b : _GEN_14728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14730 = 9'h96 == r_count_36_io_out ? io_r_150_b : _GEN_14729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14731 = 9'h97 == r_count_36_io_out ? io_r_151_b : _GEN_14730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14732 = 9'h98 == r_count_36_io_out ? io_r_152_b : _GEN_14731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14733 = 9'h99 == r_count_36_io_out ? io_r_153_b : _GEN_14732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14734 = 9'h9a == r_count_36_io_out ? io_r_154_b : _GEN_14733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14735 = 9'h9b == r_count_36_io_out ? io_r_155_b : _GEN_14734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14736 = 9'h9c == r_count_36_io_out ? io_r_156_b : _GEN_14735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14737 = 9'h9d == r_count_36_io_out ? io_r_157_b : _GEN_14736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14738 = 9'h9e == r_count_36_io_out ? io_r_158_b : _GEN_14737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14739 = 9'h9f == r_count_36_io_out ? io_r_159_b : _GEN_14738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14740 = 9'ha0 == r_count_36_io_out ? io_r_160_b : _GEN_14739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14741 = 9'ha1 == r_count_36_io_out ? io_r_161_b : _GEN_14740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14742 = 9'ha2 == r_count_36_io_out ? io_r_162_b : _GEN_14741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14743 = 9'ha3 == r_count_36_io_out ? io_r_163_b : _GEN_14742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14744 = 9'ha4 == r_count_36_io_out ? io_r_164_b : _GEN_14743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14745 = 9'ha5 == r_count_36_io_out ? io_r_165_b : _GEN_14744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14746 = 9'ha6 == r_count_36_io_out ? io_r_166_b : _GEN_14745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14747 = 9'ha7 == r_count_36_io_out ? io_r_167_b : _GEN_14746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14748 = 9'ha8 == r_count_36_io_out ? io_r_168_b : _GEN_14747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14749 = 9'ha9 == r_count_36_io_out ? io_r_169_b : _GEN_14748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14750 = 9'haa == r_count_36_io_out ? io_r_170_b : _GEN_14749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14751 = 9'hab == r_count_36_io_out ? io_r_171_b : _GEN_14750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14752 = 9'hac == r_count_36_io_out ? io_r_172_b : _GEN_14751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14753 = 9'had == r_count_36_io_out ? io_r_173_b : _GEN_14752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14754 = 9'hae == r_count_36_io_out ? io_r_174_b : _GEN_14753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14755 = 9'haf == r_count_36_io_out ? io_r_175_b : _GEN_14754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14756 = 9'hb0 == r_count_36_io_out ? io_r_176_b : _GEN_14755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14757 = 9'hb1 == r_count_36_io_out ? io_r_177_b : _GEN_14756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14758 = 9'hb2 == r_count_36_io_out ? io_r_178_b : _GEN_14757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14759 = 9'hb3 == r_count_36_io_out ? io_r_179_b : _GEN_14758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14760 = 9'hb4 == r_count_36_io_out ? io_r_180_b : _GEN_14759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14761 = 9'hb5 == r_count_36_io_out ? io_r_181_b : _GEN_14760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14762 = 9'hb6 == r_count_36_io_out ? io_r_182_b : _GEN_14761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14763 = 9'hb7 == r_count_36_io_out ? io_r_183_b : _GEN_14762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14764 = 9'hb8 == r_count_36_io_out ? io_r_184_b : _GEN_14763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14765 = 9'hb9 == r_count_36_io_out ? io_r_185_b : _GEN_14764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14766 = 9'hba == r_count_36_io_out ? io_r_186_b : _GEN_14765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14767 = 9'hbb == r_count_36_io_out ? io_r_187_b : _GEN_14766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14768 = 9'hbc == r_count_36_io_out ? io_r_188_b : _GEN_14767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14769 = 9'hbd == r_count_36_io_out ? io_r_189_b : _GEN_14768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14770 = 9'hbe == r_count_36_io_out ? io_r_190_b : _GEN_14769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14771 = 9'hbf == r_count_36_io_out ? io_r_191_b : _GEN_14770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14772 = 9'hc0 == r_count_36_io_out ? io_r_192_b : _GEN_14771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14773 = 9'hc1 == r_count_36_io_out ? io_r_193_b : _GEN_14772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14774 = 9'hc2 == r_count_36_io_out ? io_r_194_b : _GEN_14773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14775 = 9'hc3 == r_count_36_io_out ? io_r_195_b : _GEN_14774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14776 = 9'hc4 == r_count_36_io_out ? io_r_196_b : _GEN_14775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14777 = 9'hc5 == r_count_36_io_out ? io_r_197_b : _GEN_14776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14778 = 9'hc6 == r_count_36_io_out ? io_r_198_b : _GEN_14777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14779 = 9'hc7 == r_count_36_io_out ? io_r_199_b : _GEN_14778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14780 = 9'hc8 == r_count_36_io_out ? io_r_200_b : _GEN_14779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14781 = 9'hc9 == r_count_36_io_out ? io_r_201_b : _GEN_14780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14782 = 9'hca == r_count_36_io_out ? io_r_202_b : _GEN_14781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14783 = 9'hcb == r_count_36_io_out ? io_r_203_b : _GEN_14782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14784 = 9'hcc == r_count_36_io_out ? io_r_204_b : _GEN_14783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14785 = 9'hcd == r_count_36_io_out ? io_r_205_b : _GEN_14784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14786 = 9'hce == r_count_36_io_out ? io_r_206_b : _GEN_14785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14787 = 9'hcf == r_count_36_io_out ? io_r_207_b : _GEN_14786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14788 = 9'hd0 == r_count_36_io_out ? io_r_208_b : _GEN_14787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14789 = 9'hd1 == r_count_36_io_out ? io_r_209_b : _GEN_14788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14790 = 9'hd2 == r_count_36_io_out ? io_r_210_b : _GEN_14789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14791 = 9'hd3 == r_count_36_io_out ? io_r_211_b : _GEN_14790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14792 = 9'hd4 == r_count_36_io_out ? io_r_212_b : _GEN_14791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14793 = 9'hd5 == r_count_36_io_out ? io_r_213_b : _GEN_14792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14794 = 9'hd6 == r_count_36_io_out ? io_r_214_b : _GEN_14793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14795 = 9'hd7 == r_count_36_io_out ? io_r_215_b : _GEN_14794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14796 = 9'hd8 == r_count_36_io_out ? io_r_216_b : _GEN_14795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14797 = 9'hd9 == r_count_36_io_out ? io_r_217_b : _GEN_14796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14798 = 9'hda == r_count_36_io_out ? io_r_218_b : _GEN_14797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14799 = 9'hdb == r_count_36_io_out ? io_r_219_b : _GEN_14798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14800 = 9'hdc == r_count_36_io_out ? io_r_220_b : _GEN_14799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14801 = 9'hdd == r_count_36_io_out ? io_r_221_b : _GEN_14800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14802 = 9'hde == r_count_36_io_out ? io_r_222_b : _GEN_14801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14803 = 9'hdf == r_count_36_io_out ? io_r_223_b : _GEN_14802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14804 = 9'he0 == r_count_36_io_out ? io_r_224_b : _GEN_14803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14805 = 9'he1 == r_count_36_io_out ? io_r_225_b : _GEN_14804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14806 = 9'he2 == r_count_36_io_out ? io_r_226_b : _GEN_14805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14807 = 9'he3 == r_count_36_io_out ? io_r_227_b : _GEN_14806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14808 = 9'he4 == r_count_36_io_out ? io_r_228_b : _GEN_14807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14809 = 9'he5 == r_count_36_io_out ? io_r_229_b : _GEN_14808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14810 = 9'he6 == r_count_36_io_out ? io_r_230_b : _GEN_14809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14811 = 9'he7 == r_count_36_io_out ? io_r_231_b : _GEN_14810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14812 = 9'he8 == r_count_36_io_out ? io_r_232_b : _GEN_14811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14813 = 9'he9 == r_count_36_io_out ? io_r_233_b : _GEN_14812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14814 = 9'hea == r_count_36_io_out ? io_r_234_b : _GEN_14813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14815 = 9'heb == r_count_36_io_out ? io_r_235_b : _GEN_14814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14816 = 9'hec == r_count_36_io_out ? io_r_236_b : _GEN_14815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14817 = 9'hed == r_count_36_io_out ? io_r_237_b : _GEN_14816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14818 = 9'hee == r_count_36_io_out ? io_r_238_b : _GEN_14817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14819 = 9'hef == r_count_36_io_out ? io_r_239_b : _GEN_14818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14820 = 9'hf0 == r_count_36_io_out ? io_r_240_b : _GEN_14819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14821 = 9'hf1 == r_count_36_io_out ? io_r_241_b : _GEN_14820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14822 = 9'hf2 == r_count_36_io_out ? io_r_242_b : _GEN_14821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14823 = 9'hf3 == r_count_36_io_out ? io_r_243_b : _GEN_14822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14824 = 9'hf4 == r_count_36_io_out ? io_r_244_b : _GEN_14823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14825 = 9'hf5 == r_count_36_io_out ? io_r_245_b : _GEN_14824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14826 = 9'hf6 == r_count_36_io_out ? io_r_246_b : _GEN_14825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14827 = 9'hf7 == r_count_36_io_out ? io_r_247_b : _GEN_14826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14828 = 9'hf8 == r_count_36_io_out ? io_r_248_b : _GEN_14827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14829 = 9'hf9 == r_count_36_io_out ? io_r_249_b : _GEN_14828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14830 = 9'hfa == r_count_36_io_out ? io_r_250_b : _GEN_14829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14831 = 9'hfb == r_count_36_io_out ? io_r_251_b : _GEN_14830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14832 = 9'hfc == r_count_36_io_out ? io_r_252_b : _GEN_14831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14833 = 9'hfd == r_count_36_io_out ? io_r_253_b : _GEN_14832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14834 = 9'hfe == r_count_36_io_out ? io_r_254_b : _GEN_14833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14835 = 9'hff == r_count_36_io_out ? io_r_255_b : _GEN_14834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14836 = 9'h100 == r_count_36_io_out ? io_r_256_b : _GEN_14835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14837 = 9'h101 == r_count_36_io_out ? io_r_257_b : _GEN_14836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14838 = 9'h102 == r_count_36_io_out ? io_r_258_b : _GEN_14837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14839 = 9'h103 == r_count_36_io_out ? io_r_259_b : _GEN_14838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14840 = 9'h104 == r_count_36_io_out ? io_r_260_b : _GEN_14839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14841 = 9'h105 == r_count_36_io_out ? io_r_261_b : _GEN_14840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14842 = 9'h106 == r_count_36_io_out ? io_r_262_b : _GEN_14841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14843 = 9'h107 == r_count_36_io_out ? io_r_263_b : _GEN_14842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14844 = 9'h108 == r_count_36_io_out ? io_r_264_b : _GEN_14843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14845 = 9'h109 == r_count_36_io_out ? io_r_265_b : _GEN_14844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14846 = 9'h10a == r_count_36_io_out ? io_r_266_b : _GEN_14845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14847 = 9'h10b == r_count_36_io_out ? io_r_267_b : _GEN_14846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14848 = 9'h10c == r_count_36_io_out ? io_r_268_b : _GEN_14847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14849 = 9'h10d == r_count_36_io_out ? io_r_269_b : _GEN_14848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14850 = 9'h10e == r_count_36_io_out ? io_r_270_b : _GEN_14849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14851 = 9'h10f == r_count_36_io_out ? io_r_271_b : _GEN_14850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14852 = 9'h110 == r_count_36_io_out ? io_r_272_b : _GEN_14851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14853 = 9'h111 == r_count_36_io_out ? io_r_273_b : _GEN_14852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14854 = 9'h112 == r_count_36_io_out ? io_r_274_b : _GEN_14853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14855 = 9'h113 == r_count_36_io_out ? io_r_275_b : _GEN_14854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14856 = 9'h114 == r_count_36_io_out ? io_r_276_b : _GEN_14855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14857 = 9'h115 == r_count_36_io_out ? io_r_277_b : _GEN_14856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14858 = 9'h116 == r_count_36_io_out ? io_r_278_b : _GEN_14857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14859 = 9'h117 == r_count_36_io_out ? io_r_279_b : _GEN_14858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14860 = 9'h118 == r_count_36_io_out ? io_r_280_b : _GEN_14859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14861 = 9'h119 == r_count_36_io_out ? io_r_281_b : _GEN_14860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14862 = 9'h11a == r_count_36_io_out ? io_r_282_b : _GEN_14861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14863 = 9'h11b == r_count_36_io_out ? io_r_283_b : _GEN_14862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14864 = 9'h11c == r_count_36_io_out ? io_r_284_b : _GEN_14863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14865 = 9'h11d == r_count_36_io_out ? io_r_285_b : _GEN_14864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14866 = 9'h11e == r_count_36_io_out ? io_r_286_b : _GEN_14865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14867 = 9'h11f == r_count_36_io_out ? io_r_287_b : _GEN_14866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14868 = 9'h120 == r_count_36_io_out ? io_r_288_b : _GEN_14867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14869 = 9'h121 == r_count_36_io_out ? io_r_289_b : _GEN_14868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14870 = 9'h122 == r_count_36_io_out ? io_r_290_b : _GEN_14869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14871 = 9'h123 == r_count_36_io_out ? io_r_291_b : _GEN_14870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14872 = 9'h124 == r_count_36_io_out ? io_r_292_b : _GEN_14871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14873 = 9'h125 == r_count_36_io_out ? io_r_293_b : _GEN_14872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14874 = 9'h126 == r_count_36_io_out ? io_r_294_b : _GEN_14873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14875 = 9'h127 == r_count_36_io_out ? io_r_295_b : _GEN_14874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14876 = 9'h128 == r_count_36_io_out ? io_r_296_b : _GEN_14875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14877 = 9'h129 == r_count_36_io_out ? io_r_297_b : _GEN_14876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14878 = 9'h12a == r_count_36_io_out ? io_r_298_b : _GEN_14877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14879 = 9'h12b == r_count_36_io_out ? io_r_299_b : _GEN_14878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14880 = 9'h12c == r_count_36_io_out ? io_r_300_b : _GEN_14879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14881 = 9'h12d == r_count_36_io_out ? io_r_301_b : _GEN_14880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14882 = 9'h12e == r_count_36_io_out ? io_r_302_b : _GEN_14881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14883 = 9'h12f == r_count_36_io_out ? io_r_303_b : _GEN_14882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14884 = 9'h130 == r_count_36_io_out ? io_r_304_b : _GEN_14883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14885 = 9'h131 == r_count_36_io_out ? io_r_305_b : _GEN_14884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14886 = 9'h132 == r_count_36_io_out ? io_r_306_b : _GEN_14885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14887 = 9'h133 == r_count_36_io_out ? io_r_307_b : _GEN_14886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14888 = 9'h134 == r_count_36_io_out ? io_r_308_b : _GEN_14887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14889 = 9'h135 == r_count_36_io_out ? io_r_309_b : _GEN_14888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14890 = 9'h136 == r_count_36_io_out ? io_r_310_b : _GEN_14889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14891 = 9'h137 == r_count_36_io_out ? io_r_311_b : _GEN_14890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14892 = 9'h138 == r_count_36_io_out ? io_r_312_b : _GEN_14891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14893 = 9'h139 == r_count_36_io_out ? io_r_313_b : _GEN_14892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14894 = 9'h13a == r_count_36_io_out ? io_r_314_b : _GEN_14893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14895 = 9'h13b == r_count_36_io_out ? io_r_315_b : _GEN_14894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14896 = 9'h13c == r_count_36_io_out ? io_r_316_b : _GEN_14895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14897 = 9'h13d == r_count_36_io_out ? io_r_317_b : _GEN_14896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14898 = 9'h13e == r_count_36_io_out ? io_r_318_b : _GEN_14897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14899 = 9'h13f == r_count_36_io_out ? io_r_319_b : _GEN_14898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14900 = 9'h140 == r_count_36_io_out ? io_r_320_b : _GEN_14899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14901 = 9'h141 == r_count_36_io_out ? io_r_321_b : _GEN_14900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14902 = 9'h142 == r_count_36_io_out ? io_r_322_b : _GEN_14901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14903 = 9'h143 == r_count_36_io_out ? io_r_323_b : _GEN_14902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14904 = 9'h144 == r_count_36_io_out ? io_r_324_b : _GEN_14903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14905 = 9'h145 == r_count_36_io_out ? io_r_325_b : _GEN_14904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14906 = 9'h146 == r_count_36_io_out ? io_r_326_b : _GEN_14905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14907 = 9'h147 == r_count_36_io_out ? io_r_327_b : _GEN_14906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14908 = 9'h148 == r_count_36_io_out ? io_r_328_b : _GEN_14907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14909 = 9'h149 == r_count_36_io_out ? io_r_329_b : _GEN_14908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14910 = 9'h14a == r_count_36_io_out ? io_r_330_b : _GEN_14909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14911 = 9'h14b == r_count_36_io_out ? io_r_331_b : _GEN_14910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14912 = 9'h14c == r_count_36_io_out ? io_r_332_b : _GEN_14911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14913 = 9'h14d == r_count_36_io_out ? io_r_333_b : _GEN_14912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14914 = 9'h14e == r_count_36_io_out ? io_r_334_b : _GEN_14913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14915 = 9'h14f == r_count_36_io_out ? io_r_335_b : _GEN_14914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14916 = 9'h150 == r_count_36_io_out ? io_r_336_b : _GEN_14915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14917 = 9'h151 == r_count_36_io_out ? io_r_337_b : _GEN_14916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14918 = 9'h152 == r_count_36_io_out ? io_r_338_b : _GEN_14917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14919 = 9'h153 == r_count_36_io_out ? io_r_339_b : _GEN_14918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14920 = 9'h154 == r_count_36_io_out ? io_r_340_b : _GEN_14919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14921 = 9'h155 == r_count_36_io_out ? io_r_341_b : _GEN_14920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14922 = 9'h156 == r_count_36_io_out ? io_r_342_b : _GEN_14921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14923 = 9'h157 == r_count_36_io_out ? io_r_343_b : _GEN_14922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14924 = 9'h158 == r_count_36_io_out ? io_r_344_b : _GEN_14923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14925 = 9'h159 == r_count_36_io_out ? io_r_345_b : _GEN_14924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14926 = 9'h15a == r_count_36_io_out ? io_r_346_b : _GEN_14925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14927 = 9'h15b == r_count_36_io_out ? io_r_347_b : _GEN_14926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14928 = 9'h15c == r_count_36_io_out ? io_r_348_b : _GEN_14927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14929 = 9'h15d == r_count_36_io_out ? io_r_349_b : _GEN_14928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14930 = 9'h15e == r_count_36_io_out ? io_r_350_b : _GEN_14929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14931 = 9'h15f == r_count_36_io_out ? io_r_351_b : _GEN_14930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14932 = 9'h160 == r_count_36_io_out ? io_r_352_b : _GEN_14931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14933 = 9'h161 == r_count_36_io_out ? io_r_353_b : _GEN_14932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14934 = 9'h162 == r_count_36_io_out ? io_r_354_b : _GEN_14933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14935 = 9'h163 == r_count_36_io_out ? io_r_355_b : _GEN_14934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14936 = 9'h164 == r_count_36_io_out ? io_r_356_b : _GEN_14935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14937 = 9'h165 == r_count_36_io_out ? io_r_357_b : _GEN_14936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14938 = 9'h166 == r_count_36_io_out ? io_r_358_b : _GEN_14937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14939 = 9'h167 == r_count_36_io_out ? io_r_359_b : _GEN_14938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14940 = 9'h168 == r_count_36_io_out ? io_r_360_b : _GEN_14939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14941 = 9'h169 == r_count_36_io_out ? io_r_361_b : _GEN_14940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14942 = 9'h16a == r_count_36_io_out ? io_r_362_b : _GEN_14941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14943 = 9'h16b == r_count_36_io_out ? io_r_363_b : _GEN_14942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14944 = 9'h16c == r_count_36_io_out ? io_r_364_b : _GEN_14943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14945 = 9'h16d == r_count_36_io_out ? io_r_365_b : _GEN_14944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14946 = 9'h16e == r_count_36_io_out ? io_r_366_b : _GEN_14945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14947 = 9'h16f == r_count_36_io_out ? io_r_367_b : _GEN_14946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14948 = 9'h170 == r_count_36_io_out ? io_r_368_b : _GEN_14947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14949 = 9'h171 == r_count_36_io_out ? io_r_369_b : _GEN_14948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14950 = 9'h172 == r_count_36_io_out ? io_r_370_b : _GEN_14949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14951 = 9'h173 == r_count_36_io_out ? io_r_371_b : _GEN_14950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14952 = 9'h174 == r_count_36_io_out ? io_r_372_b : _GEN_14951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14953 = 9'h175 == r_count_36_io_out ? io_r_373_b : _GEN_14952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14954 = 9'h176 == r_count_36_io_out ? io_r_374_b : _GEN_14953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14955 = 9'h177 == r_count_36_io_out ? io_r_375_b : _GEN_14954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14956 = 9'h178 == r_count_36_io_out ? io_r_376_b : _GEN_14955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14957 = 9'h179 == r_count_36_io_out ? io_r_377_b : _GEN_14956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14958 = 9'h17a == r_count_36_io_out ? io_r_378_b : _GEN_14957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14959 = 9'h17b == r_count_36_io_out ? io_r_379_b : _GEN_14958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14960 = 9'h17c == r_count_36_io_out ? io_r_380_b : _GEN_14959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14961 = 9'h17d == r_count_36_io_out ? io_r_381_b : _GEN_14960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14962 = 9'h17e == r_count_36_io_out ? io_r_382_b : _GEN_14961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14963 = 9'h17f == r_count_36_io_out ? io_r_383_b : _GEN_14962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14964 = 9'h180 == r_count_36_io_out ? io_r_384_b : _GEN_14963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14965 = 9'h181 == r_count_36_io_out ? io_r_385_b : _GEN_14964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14966 = 9'h182 == r_count_36_io_out ? io_r_386_b : _GEN_14965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14967 = 9'h183 == r_count_36_io_out ? io_r_387_b : _GEN_14966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14968 = 9'h184 == r_count_36_io_out ? io_r_388_b : _GEN_14967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14969 = 9'h185 == r_count_36_io_out ? io_r_389_b : _GEN_14968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14970 = 9'h186 == r_count_36_io_out ? io_r_390_b : _GEN_14969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14971 = 9'h187 == r_count_36_io_out ? io_r_391_b : _GEN_14970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14972 = 9'h188 == r_count_36_io_out ? io_r_392_b : _GEN_14971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14973 = 9'h189 == r_count_36_io_out ? io_r_393_b : _GEN_14972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14974 = 9'h18a == r_count_36_io_out ? io_r_394_b : _GEN_14973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14975 = 9'h18b == r_count_36_io_out ? io_r_395_b : _GEN_14974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14976 = 9'h18c == r_count_36_io_out ? io_r_396_b : _GEN_14975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14977 = 9'h18d == r_count_36_io_out ? io_r_397_b : _GEN_14976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14978 = 9'h18e == r_count_36_io_out ? io_r_398_b : _GEN_14977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14981 = 9'h1 == r_count_37_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14982 = 9'h2 == r_count_37_io_out ? io_r_2_b : _GEN_14981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14983 = 9'h3 == r_count_37_io_out ? io_r_3_b : _GEN_14982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14984 = 9'h4 == r_count_37_io_out ? io_r_4_b : _GEN_14983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14985 = 9'h5 == r_count_37_io_out ? io_r_5_b : _GEN_14984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14986 = 9'h6 == r_count_37_io_out ? io_r_6_b : _GEN_14985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14987 = 9'h7 == r_count_37_io_out ? io_r_7_b : _GEN_14986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14988 = 9'h8 == r_count_37_io_out ? io_r_8_b : _GEN_14987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14989 = 9'h9 == r_count_37_io_out ? io_r_9_b : _GEN_14988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14990 = 9'ha == r_count_37_io_out ? io_r_10_b : _GEN_14989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14991 = 9'hb == r_count_37_io_out ? io_r_11_b : _GEN_14990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14992 = 9'hc == r_count_37_io_out ? io_r_12_b : _GEN_14991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14993 = 9'hd == r_count_37_io_out ? io_r_13_b : _GEN_14992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14994 = 9'he == r_count_37_io_out ? io_r_14_b : _GEN_14993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14995 = 9'hf == r_count_37_io_out ? io_r_15_b : _GEN_14994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14996 = 9'h10 == r_count_37_io_out ? io_r_16_b : _GEN_14995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14997 = 9'h11 == r_count_37_io_out ? io_r_17_b : _GEN_14996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14998 = 9'h12 == r_count_37_io_out ? io_r_18_b : _GEN_14997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14999 = 9'h13 == r_count_37_io_out ? io_r_19_b : _GEN_14998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15000 = 9'h14 == r_count_37_io_out ? io_r_20_b : _GEN_14999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15001 = 9'h15 == r_count_37_io_out ? io_r_21_b : _GEN_15000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15002 = 9'h16 == r_count_37_io_out ? io_r_22_b : _GEN_15001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15003 = 9'h17 == r_count_37_io_out ? io_r_23_b : _GEN_15002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15004 = 9'h18 == r_count_37_io_out ? io_r_24_b : _GEN_15003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15005 = 9'h19 == r_count_37_io_out ? io_r_25_b : _GEN_15004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15006 = 9'h1a == r_count_37_io_out ? io_r_26_b : _GEN_15005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15007 = 9'h1b == r_count_37_io_out ? io_r_27_b : _GEN_15006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15008 = 9'h1c == r_count_37_io_out ? io_r_28_b : _GEN_15007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15009 = 9'h1d == r_count_37_io_out ? io_r_29_b : _GEN_15008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15010 = 9'h1e == r_count_37_io_out ? io_r_30_b : _GEN_15009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15011 = 9'h1f == r_count_37_io_out ? io_r_31_b : _GEN_15010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15012 = 9'h20 == r_count_37_io_out ? io_r_32_b : _GEN_15011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15013 = 9'h21 == r_count_37_io_out ? io_r_33_b : _GEN_15012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15014 = 9'h22 == r_count_37_io_out ? io_r_34_b : _GEN_15013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15015 = 9'h23 == r_count_37_io_out ? io_r_35_b : _GEN_15014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15016 = 9'h24 == r_count_37_io_out ? io_r_36_b : _GEN_15015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15017 = 9'h25 == r_count_37_io_out ? io_r_37_b : _GEN_15016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15018 = 9'h26 == r_count_37_io_out ? io_r_38_b : _GEN_15017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15019 = 9'h27 == r_count_37_io_out ? io_r_39_b : _GEN_15018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15020 = 9'h28 == r_count_37_io_out ? io_r_40_b : _GEN_15019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15021 = 9'h29 == r_count_37_io_out ? io_r_41_b : _GEN_15020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15022 = 9'h2a == r_count_37_io_out ? io_r_42_b : _GEN_15021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15023 = 9'h2b == r_count_37_io_out ? io_r_43_b : _GEN_15022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15024 = 9'h2c == r_count_37_io_out ? io_r_44_b : _GEN_15023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15025 = 9'h2d == r_count_37_io_out ? io_r_45_b : _GEN_15024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15026 = 9'h2e == r_count_37_io_out ? io_r_46_b : _GEN_15025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15027 = 9'h2f == r_count_37_io_out ? io_r_47_b : _GEN_15026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15028 = 9'h30 == r_count_37_io_out ? io_r_48_b : _GEN_15027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15029 = 9'h31 == r_count_37_io_out ? io_r_49_b : _GEN_15028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15030 = 9'h32 == r_count_37_io_out ? io_r_50_b : _GEN_15029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15031 = 9'h33 == r_count_37_io_out ? io_r_51_b : _GEN_15030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15032 = 9'h34 == r_count_37_io_out ? io_r_52_b : _GEN_15031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15033 = 9'h35 == r_count_37_io_out ? io_r_53_b : _GEN_15032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15034 = 9'h36 == r_count_37_io_out ? io_r_54_b : _GEN_15033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15035 = 9'h37 == r_count_37_io_out ? io_r_55_b : _GEN_15034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15036 = 9'h38 == r_count_37_io_out ? io_r_56_b : _GEN_15035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15037 = 9'h39 == r_count_37_io_out ? io_r_57_b : _GEN_15036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15038 = 9'h3a == r_count_37_io_out ? io_r_58_b : _GEN_15037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15039 = 9'h3b == r_count_37_io_out ? io_r_59_b : _GEN_15038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15040 = 9'h3c == r_count_37_io_out ? io_r_60_b : _GEN_15039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15041 = 9'h3d == r_count_37_io_out ? io_r_61_b : _GEN_15040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15042 = 9'h3e == r_count_37_io_out ? io_r_62_b : _GEN_15041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15043 = 9'h3f == r_count_37_io_out ? io_r_63_b : _GEN_15042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15044 = 9'h40 == r_count_37_io_out ? io_r_64_b : _GEN_15043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15045 = 9'h41 == r_count_37_io_out ? io_r_65_b : _GEN_15044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15046 = 9'h42 == r_count_37_io_out ? io_r_66_b : _GEN_15045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15047 = 9'h43 == r_count_37_io_out ? io_r_67_b : _GEN_15046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15048 = 9'h44 == r_count_37_io_out ? io_r_68_b : _GEN_15047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15049 = 9'h45 == r_count_37_io_out ? io_r_69_b : _GEN_15048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15050 = 9'h46 == r_count_37_io_out ? io_r_70_b : _GEN_15049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15051 = 9'h47 == r_count_37_io_out ? io_r_71_b : _GEN_15050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15052 = 9'h48 == r_count_37_io_out ? io_r_72_b : _GEN_15051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15053 = 9'h49 == r_count_37_io_out ? io_r_73_b : _GEN_15052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15054 = 9'h4a == r_count_37_io_out ? io_r_74_b : _GEN_15053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15055 = 9'h4b == r_count_37_io_out ? io_r_75_b : _GEN_15054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15056 = 9'h4c == r_count_37_io_out ? io_r_76_b : _GEN_15055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15057 = 9'h4d == r_count_37_io_out ? io_r_77_b : _GEN_15056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15058 = 9'h4e == r_count_37_io_out ? io_r_78_b : _GEN_15057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15059 = 9'h4f == r_count_37_io_out ? io_r_79_b : _GEN_15058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15060 = 9'h50 == r_count_37_io_out ? io_r_80_b : _GEN_15059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15061 = 9'h51 == r_count_37_io_out ? io_r_81_b : _GEN_15060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15062 = 9'h52 == r_count_37_io_out ? io_r_82_b : _GEN_15061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15063 = 9'h53 == r_count_37_io_out ? io_r_83_b : _GEN_15062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15064 = 9'h54 == r_count_37_io_out ? io_r_84_b : _GEN_15063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15065 = 9'h55 == r_count_37_io_out ? io_r_85_b : _GEN_15064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15066 = 9'h56 == r_count_37_io_out ? io_r_86_b : _GEN_15065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15067 = 9'h57 == r_count_37_io_out ? io_r_87_b : _GEN_15066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15068 = 9'h58 == r_count_37_io_out ? io_r_88_b : _GEN_15067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15069 = 9'h59 == r_count_37_io_out ? io_r_89_b : _GEN_15068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15070 = 9'h5a == r_count_37_io_out ? io_r_90_b : _GEN_15069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15071 = 9'h5b == r_count_37_io_out ? io_r_91_b : _GEN_15070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15072 = 9'h5c == r_count_37_io_out ? io_r_92_b : _GEN_15071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15073 = 9'h5d == r_count_37_io_out ? io_r_93_b : _GEN_15072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15074 = 9'h5e == r_count_37_io_out ? io_r_94_b : _GEN_15073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15075 = 9'h5f == r_count_37_io_out ? io_r_95_b : _GEN_15074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15076 = 9'h60 == r_count_37_io_out ? io_r_96_b : _GEN_15075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15077 = 9'h61 == r_count_37_io_out ? io_r_97_b : _GEN_15076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15078 = 9'h62 == r_count_37_io_out ? io_r_98_b : _GEN_15077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15079 = 9'h63 == r_count_37_io_out ? io_r_99_b : _GEN_15078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15080 = 9'h64 == r_count_37_io_out ? io_r_100_b : _GEN_15079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15081 = 9'h65 == r_count_37_io_out ? io_r_101_b : _GEN_15080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15082 = 9'h66 == r_count_37_io_out ? io_r_102_b : _GEN_15081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15083 = 9'h67 == r_count_37_io_out ? io_r_103_b : _GEN_15082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15084 = 9'h68 == r_count_37_io_out ? io_r_104_b : _GEN_15083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15085 = 9'h69 == r_count_37_io_out ? io_r_105_b : _GEN_15084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15086 = 9'h6a == r_count_37_io_out ? io_r_106_b : _GEN_15085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15087 = 9'h6b == r_count_37_io_out ? io_r_107_b : _GEN_15086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15088 = 9'h6c == r_count_37_io_out ? io_r_108_b : _GEN_15087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15089 = 9'h6d == r_count_37_io_out ? io_r_109_b : _GEN_15088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15090 = 9'h6e == r_count_37_io_out ? io_r_110_b : _GEN_15089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15091 = 9'h6f == r_count_37_io_out ? io_r_111_b : _GEN_15090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15092 = 9'h70 == r_count_37_io_out ? io_r_112_b : _GEN_15091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15093 = 9'h71 == r_count_37_io_out ? io_r_113_b : _GEN_15092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15094 = 9'h72 == r_count_37_io_out ? io_r_114_b : _GEN_15093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15095 = 9'h73 == r_count_37_io_out ? io_r_115_b : _GEN_15094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15096 = 9'h74 == r_count_37_io_out ? io_r_116_b : _GEN_15095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15097 = 9'h75 == r_count_37_io_out ? io_r_117_b : _GEN_15096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15098 = 9'h76 == r_count_37_io_out ? io_r_118_b : _GEN_15097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15099 = 9'h77 == r_count_37_io_out ? io_r_119_b : _GEN_15098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15100 = 9'h78 == r_count_37_io_out ? io_r_120_b : _GEN_15099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15101 = 9'h79 == r_count_37_io_out ? io_r_121_b : _GEN_15100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15102 = 9'h7a == r_count_37_io_out ? io_r_122_b : _GEN_15101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15103 = 9'h7b == r_count_37_io_out ? io_r_123_b : _GEN_15102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15104 = 9'h7c == r_count_37_io_out ? io_r_124_b : _GEN_15103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15105 = 9'h7d == r_count_37_io_out ? io_r_125_b : _GEN_15104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15106 = 9'h7e == r_count_37_io_out ? io_r_126_b : _GEN_15105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15107 = 9'h7f == r_count_37_io_out ? io_r_127_b : _GEN_15106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15108 = 9'h80 == r_count_37_io_out ? io_r_128_b : _GEN_15107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15109 = 9'h81 == r_count_37_io_out ? io_r_129_b : _GEN_15108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15110 = 9'h82 == r_count_37_io_out ? io_r_130_b : _GEN_15109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15111 = 9'h83 == r_count_37_io_out ? io_r_131_b : _GEN_15110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15112 = 9'h84 == r_count_37_io_out ? io_r_132_b : _GEN_15111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15113 = 9'h85 == r_count_37_io_out ? io_r_133_b : _GEN_15112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15114 = 9'h86 == r_count_37_io_out ? io_r_134_b : _GEN_15113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15115 = 9'h87 == r_count_37_io_out ? io_r_135_b : _GEN_15114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15116 = 9'h88 == r_count_37_io_out ? io_r_136_b : _GEN_15115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15117 = 9'h89 == r_count_37_io_out ? io_r_137_b : _GEN_15116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15118 = 9'h8a == r_count_37_io_out ? io_r_138_b : _GEN_15117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15119 = 9'h8b == r_count_37_io_out ? io_r_139_b : _GEN_15118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15120 = 9'h8c == r_count_37_io_out ? io_r_140_b : _GEN_15119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15121 = 9'h8d == r_count_37_io_out ? io_r_141_b : _GEN_15120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15122 = 9'h8e == r_count_37_io_out ? io_r_142_b : _GEN_15121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15123 = 9'h8f == r_count_37_io_out ? io_r_143_b : _GEN_15122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15124 = 9'h90 == r_count_37_io_out ? io_r_144_b : _GEN_15123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15125 = 9'h91 == r_count_37_io_out ? io_r_145_b : _GEN_15124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15126 = 9'h92 == r_count_37_io_out ? io_r_146_b : _GEN_15125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15127 = 9'h93 == r_count_37_io_out ? io_r_147_b : _GEN_15126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15128 = 9'h94 == r_count_37_io_out ? io_r_148_b : _GEN_15127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15129 = 9'h95 == r_count_37_io_out ? io_r_149_b : _GEN_15128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15130 = 9'h96 == r_count_37_io_out ? io_r_150_b : _GEN_15129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15131 = 9'h97 == r_count_37_io_out ? io_r_151_b : _GEN_15130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15132 = 9'h98 == r_count_37_io_out ? io_r_152_b : _GEN_15131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15133 = 9'h99 == r_count_37_io_out ? io_r_153_b : _GEN_15132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15134 = 9'h9a == r_count_37_io_out ? io_r_154_b : _GEN_15133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15135 = 9'h9b == r_count_37_io_out ? io_r_155_b : _GEN_15134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15136 = 9'h9c == r_count_37_io_out ? io_r_156_b : _GEN_15135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15137 = 9'h9d == r_count_37_io_out ? io_r_157_b : _GEN_15136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15138 = 9'h9e == r_count_37_io_out ? io_r_158_b : _GEN_15137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15139 = 9'h9f == r_count_37_io_out ? io_r_159_b : _GEN_15138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15140 = 9'ha0 == r_count_37_io_out ? io_r_160_b : _GEN_15139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15141 = 9'ha1 == r_count_37_io_out ? io_r_161_b : _GEN_15140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15142 = 9'ha2 == r_count_37_io_out ? io_r_162_b : _GEN_15141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15143 = 9'ha3 == r_count_37_io_out ? io_r_163_b : _GEN_15142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15144 = 9'ha4 == r_count_37_io_out ? io_r_164_b : _GEN_15143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15145 = 9'ha5 == r_count_37_io_out ? io_r_165_b : _GEN_15144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15146 = 9'ha6 == r_count_37_io_out ? io_r_166_b : _GEN_15145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15147 = 9'ha7 == r_count_37_io_out ? io_r_167_b : _GEN_15146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15148 = 9'ha8 == r_count_37_io_out ? io_r_168_b : _GEN_15147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15149 = 9'ha9 == r_count_37_io_out ? io_r_169_b : _GEN_15148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15150 = 9'haa == r_count_37_io_out ? io_r_170_b : _GEN_15149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15151 = 9'hab == r_count_37_io_out ? io_r_171_b : _GEN_15150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15152 = 9'hac == r_count_37_io_out ? io_r_172_b : _GEN_15151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15153 = 9'had == r_count_37_io_out ? io_r_173_b : _GEN_15152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15154 = 9'hae == r_count_37_io_out ? io_r_174_b : _GEN_15153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15155 = 9'haf == r_count_37_io_out ? io_r_175_b : _GEN_15154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15156 = 9'hb0 == r_count_37_io_out ? io_r_176_b : _GEN_15155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15157 = 9'hb1 == r_count_37_io_out ? io_r_177_b : _GEN_15156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15158 = 9'hb2 == r_count_37_io_out ? io_r_178_b : _GEN_15157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15159 = 9'hb3 == r_count_37_io_out ? io_r_179_b : _GEN_15158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15160 = 9'hb4 == r_count_37_io_out ? io_r_180_b : _GEN_15159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15161 = 9'hb5 == r_count_37_io_out ? io_r_181_b : _GEN_15160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15162 = 9'hb6 == r_count_37_io_out ? io_r_182_b : _GEN_15161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15163 = 9'hb7 == r_count_37_io_out ? io_r_183_b : _GEN_15162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15164 = 9'hb8 == r_count_37_io_out ? io_r_184_b : _GEN_15163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15165 = 9'hb9 == r_count_37_io_out ? io_r_185_b : _GEN_15164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15166 = 9'hba == r_count_37_io_out ? io_r_186_b : _GEN_15165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15167 = 9'hbb == r_count_37_io_out ? io_r_187_b : _GEN_15166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15168 = 9'hbc == r_count_37_io_out ? io_r_188_b : _GEN_15167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15169 = 9'hbd == r_count_37_io_out ? io_r_189_b : _GEN_15168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15170 = 9'hbe == r_count_37_io_out ? io_r_190_b : _GEN_15169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15171 = 9'hbf == r_count_37_io_out ? io_r_191_b : _GEN_15170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15172 = 9'hc0 == r_count_37_io_out ? io_r_192_b : _GEN_15171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15173 = 9'hc1 == r_count_37_io_out ? io_r_193_b : _GEN_15172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15174 = 9'hc2 == r_count_37_io_out ? io_r_194_b : _GEN_15173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15175 = 9'hc3 == r_count_37_io_out ? io_r_195_b : _GEN_15174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15176 = 9'hc4 == r_count_37_io_out ? io_r_196_b : _GEN_15175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15177 = 9'hc5 == r_count_37_io_out ? io_r_197_b : _GEN_15176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15178 = 9'hc6 == r_count_37_io_out ? io_r_198_b : _GEN_15177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15179 = 9'hc7 == r_count_37_io_out ? io_r_199_b : _GEN_15178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15180 = 9'hc8 == r_count_37_io_out ? io_r_200_b : _GEN_15179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15181 = 9'hc9 == r_count_37_io_out ? io_r_201_b : _GEN_15180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15182 = 9'hca == r_count_37_io_out ? io_r_202_b : _GEN_15181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15183 = 9'hcb == r_count_37_io_out ? io_r_203_b : _GEN_15182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15184 = 9'hcc == r_count_37_io_out ? io_r_204_b : _GEN_15183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15185 = 9'hcd == r_count_37_io_out ? io_r_205_b : _GEN_15184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15186 = 9'hce == r_count_37_io_out ? io_r_206_b : _GEN_15185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15187 = 9'hcf == r_count_37_io_out ? io_r_207_b : _GEN_15186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15188 = 9'hd0 == r_count_37_io_out ? io_r_208_b : _GEN_15187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15189 = 9'hd1 == r_count_37_io_out ? io_r_209_b : _GEN_15188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15190 = 9'hd2 == r_count_37_io_out ? io_r_210_b : _GEN_15189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15191 = 9'hd3 == r_count_37_io_out ? io_r_211_b : _GEN_15190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15192 = 9'hd4 == r_count_37_io_out ? io_r_212_b : _GEN_15191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15193 = 9'hd5 == r_count_37_io_out ? io_r_213_b : _GEN_15192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15194 = 9'hd6 == r_count_37_io_out ? io_r_214_b : _GEN_15193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15195 = 9'hd7 == r_count_37_io_out ? io_r_215_b : _GEN_15194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15196 = 9'hd8 == r_count_37_io_out ? io_r_216_b : _GEN_15195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15197 = 9'hd9 == r_count_37_io_out ? io_r_217_b : _GEN_15196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15198 = 9'hda == r_count_37_io_out ? io_r_218_b : _GEN_15197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15199 = 9'hdb == r_count_37_io_out ? io_r_219_b : _GEN_15198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15200 = 9'hdc == r_count_37_io_out ? io_r_220_b : _GEN_15199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15201 = 9'hdd == r_count_37_io_out ? io_r_221_b : _GEN_15200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15202 = 9'hde == r_count_37_io_out ? io_r_222_b : _GEN_15201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15203 = 9'hdf == r_count_37_io_out ? io_r_223_b : _GEN_15202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15204 = 9'he0 == r_count_37_io_out ? io_r_224_b : _GEN_15203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15205 = 9'he1 == r_count_37_io_out ? io_r_225_b : _GEN_15204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15206 = 9'he2 == r_count_37_io_out ? io_r_226_b : _GEN_15205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15207 = 9'he3 == r_count_37_io_out ? io_r_227_b : _GEN_15206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15208 = 9'he4 == r_count_37_io_out ? io_r_228_b : _GEN_15207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15209 = 9'he5 == r_count_37_io_out ? io_r_229_b : _GEN_15208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15210 = 9'he6 == r_count_37_io_out ? io_r_230_b : _GEN_15209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15211 = 9'he7 == r_count_37_io_out ? io_r_231_b : _GEN_15210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15212 = 9'he8 == r_count_37_io_out ? io_r_232_b : _GEN_15211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15213 = 9'he9 == r_count_37_io_out ? io_r_233_b : _GEN_15212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15214 = 9'hea == r_count_37_io_out ? io_r_234_b : _GEN_15213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15215 = 9'heb == r_count_37_io_out ? io_r_235_b : _GEN_15214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15216 = 9'hec == r_count_37_io_out ? io_r_236_b : _GEN_15215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15217 = 9'hed == r_count_37_io_out ? io_r_237_b : _GEN_15216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15218 = 9'hee == r_count_37_io_out ? io_r_238_b : _GEN_15217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15219 = 9'hef == r_count_37_io_out ? io_r_239_b : _GEN_15218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15220 = 9'hf0 == r_count_37_io_out ? io_r_240_b : _GEN_15219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15221 = 9'hf1 == r_count_37_io_out ? io_r_241_b : _GEN_15220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15222 = 9'hf2 == r_count_37_io_out ? io_r_242_b : _GEN_15221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15223 = 9'hf3 == r_count_37_io_out ? io_r_243_b : _GEN_15222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15224 = 9'hf4 == r_count_37_io_out ? io_r_244_b : _GEN_15223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15225 = 9'hf5 == r_count_37_io_out ? io_r_245_b : _GEN_15224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15226 = 9'hf6 == r_count_37_io_out ? io_r_246_b : _GEN_15225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15227 = 9'hf7 == r_count_37_io_out ? io_r_247_b : _GEN_15226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15228 = 9'hf8 == r_count_37_io_out ? io_r_248_b : _GEN_15227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15229 = 9'hf9 == r_count_37_io_out ? io_r_249_b : _GEN_15228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15230 = 9'hfa == r_count_37_io_out ? io_r_250_b : _GEN_15229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15231 = 9'hfb == r_count_37_io_out ? io_r_251_b : _GEN_15230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15232 = 9'hfc == r_count_37_io_out ? io_r_252_b : _GEN_15231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15233 = 9'hfd == r_count_37_io_out ? io_r_253_b : _GEN_15232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15234 = 9'hfe == r_count_37_io_out ? io_r_254_b : _GEN_15233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15235 = 9'hff == r_count_37_io_out ? io_r_255_b : _GEN_15234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15236 = 9'h100 == r_count_37_io_out ? io_r_256_b : _GEN_15235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15237 = 9'h101 == r_count_37_io_out ? io_r_257_b : _GEN_15236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15238 = 9'h102 == r_count_37_io_out ? io_r_258_b : _GEN_15237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15239 = 9'h103 == r_count_37_io_out ? io_r_259_b : _GEN_15238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15240 = 9'h104 == r_count_37_io_out ? io_r_260_b : _GEN_15239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15241 = 9'h105 == r_count_37_io_out ? io_r_261_b : _GEN_15240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15242 = 9'h106 == r_count_37_io_out ? io_r_262_b : _GEN_15241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15243 = 9'h107 == r_count_37_io_out ? io_r_263_b : _GEN_15242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15244 = 9'h108 == r_count_37_io_out ? io_r_264_b : _GEN_15243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15245 = 9'h109 == r_count_37_io_out ? io_r_265_b : _GEN_15244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15246 = 9'h10a == r_count_37_io_out ? io_r_266_b : _GEN_15245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15247 = 9'h10b == r_count_37_io_out ? io_r_267_b : _GEN_15246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15248 = 9'h10c == r_count_37_io_out ? io_r_268_b : _GEN_15247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15249 = 9'h10d == r_count_37_io_out ? io_r_269_b : _GEN_15248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15250 = 9'h10e == r_count_37_io_out ? io_r_270_b : _GEN_15249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15251 = 9'h10f == r_count_37_io_out ? io_r_271_b : _GEN_15250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15252 = 9'h110 == r_count_37_io_out ? io_r_272_b : _GEN_15251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15253 = 9'h111 == r_count_37_io_out ? io_r_273_b : _GEN_15252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15254 = 9'h112 == r_count_37_io_out ? io_r_274_b : _GEN_15253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15255 = 9'h113 == r_count_37_io_out ? io_r_275_b : _GEN_15254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15256 = 9'h114 == r_count_37_io_out ? io_r_276_b : _GEN_15255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15257 = 9'h115 == r_count_37_io_out ? io_r_277_b : _GEN_15256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15258 = 9'h116 == r_count_37_io_out ? io_r_278_b : _GEN_15257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15259 = 9'h117 == r_count_37_io_out ? io_r_279_b : _GEN_15258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15260 = 9'h118 == r_count_37_io_out ? io_r_280_b : _GEN_15259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15261 = 9'h119 == r_count_37_io_out ? io_r_281_b : _GEN_15260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15262 = 9'h11a == r_count_37_io_out ? io_r_282_b : _GEN_15261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15263 = 9'h11b == r_count_37_io_out ? io_r_283_b : _GEN_15262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15264 = 9'h11c == r_count_37_io_out ? io_r_284_b : _GEN_15263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15265 = 9'h11d == r_count_37_io_out ? io_r_285_b : _GEN_15264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15266 = 9'h11e == r_count_37_io_out ? io_r_286_b : _GEN_15265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15267 = 9'h11f == r_count_37_io_out ? io_r_287_b : _GEN_15266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15268 = 9'h120 == r_count_37_io_out ? io_r_288_b : _GEN_15267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15269 = 9'h121 == r_count_37_io_out ? io_r_289_b : _GEN_15268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15270 = 9'h122 == r_count_37_io_out ? io_r_290_b : _GEN_15269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15271 = 9'h123 == r_count_37_io_out ? io_r_291_b : _GEN_15270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15272 = 9'h124 == r_count_37_io_out ? io_r_292_b : _GEN_15271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15273 = 9'h125 == r_count_37_io_out ? io_r_293_b : _GEN_15272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15274 = 9'h126 == r_count_37_io_out ? io_r_294_b : _GEN_15273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15275 = 9'h127 == r_count_37_io_out ? io_r_295_b : _GEN_15274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15276 = 9'h128 == r_count_37_io_out ? io_r_296_b : _GEN_15275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15277 = 9'h129 == r_count_37_io_out ? io_r_297_b : _GEN_15276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15278 = 9'h12a == r_count_37_io_out ? io_r_298_b : _GEN_15277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15279 = 9'h12b == r_count_37_io_out ? io_r_299_b : _GEN_15278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15280 = 9'h12c == r_count_37_io_out ? io_r_300_b : _GEN_15279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15281 = 9'h12d == r_count_37_io_out ? io_r_301_b : _GEN_15280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15282 = 9'h12e == r_count_37_io_out ? io_r_302_b : _GEN_15281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15283 = 9'h12f == r_count_37_io_out ? io_r_303_b : _GEN_15282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15284 = 9'h130 == r_count_37_io_out ? io_r_304_b : _GEN_15283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15285 = 9'h131 == r_count_37_io_out ? io_r_305_b : _GEN_15284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15286 = 9'h132 == r_count_37_io_out ? io_r_306_b : _GEN_15285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15287 = 9'h133 == r_count_37_io_out ? io_r_307_b : _GEN_15286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15288 = 9'h134 == r_count_37_io_out ? io_r_308_b : _GEN_15287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15289 = 9'h135 == r_count_37_io_out ? io_r_309_b : _GEN_15288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15290 = 9'h136 == r_count_37_io_out ? io_r_310_b : _GEN_15289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15291 = 9'h137 == r_count_37_io_out ? io_r_311_b : _GEN_15290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15292 = 9'h138 == r_count_37_io_out ? io_r_312_b : _GEN_15291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15293 = 9'h139 == r_count_37_io_out ? io_r_313_b : _GEN_15292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15294 = 9'h13a == r_count_37_io_out ? io_r_314_b : _GEN_15293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15295 = 9'h13b == r_count_37_io_out ? io_r_315_b : _GEN_15294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15296 = 9'h13c == r_count_37_io_out ? io_r_316_b : _GEN_15295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15297 = 9'h13d == r_count_37_io_out ? io_r_317_b : _GEN_15296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15298 = 9'h13e == r_count_37_io_out ? io_r_318_b : _GEN_15297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15299 = 9'h13f == r_count_37_io_out ? io_r_319_b : _GEN_15298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15300 = 9'h140 == r_count_37_io_out ? io_r_320_b : _GEN_15299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15301 = 9'h141 == r_count_37_io_out ? io_r_321_b : _GEN_15300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15302 = 9'h142 == r_count_37_io_out ? io_r_322_b : _GEN_15301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15303 = 9'h143 == r_count_37_io_out ? io_r_323_b : _GEN_15302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15304 = 9'h144 == r_count_37_io_out ? io_r_324_b : _GEN_15303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15305 = 9'h145 == r_count_37_io_out ? io_r_325_b : _GEN_15304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15306 = 9'h146 == r_count_37_io_out ? io_r_326_b : _GEN_15305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15307 = 9'h147 == r_count_37_io_out ? io_r_327_b : _GEN_15306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15308 = 9'h148 == r_count_37_io_out ? io_r_328_b : _GEN_15307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15309 = 9'h149 == r_count_37_io_out ? io_r_329_b : _GEN_15308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15310 = 9'h14a == r_count_37_io_out ? io_r_330_b : _GEN_15309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15311 = 9'h14b == r_count_37_io_out ? io_r_331_b : _GEN_15310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15312 = 9'h14c == r_count_37_io_out ? io_r_332_b : _GEN_15311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15313 = 9'h14d == r_count_37_io_out ? io_r_333_b : _GEN_15312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15314 = 9'h14e == r_count_37_io_out ? io_r_334_b : _GEN_15313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15315 = 9'h14f == r_count_37_io_out ? io_r_335_b : _GEN_15314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15316 = 9'h150 == r_count_37_io_out ? io_r_336_b : _GEN_15315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15317 = 9'h151 == r_count_37_io_out ? io_r_337_b : _GEN_15316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15318 = 9'h152 == r_count_37_io_out ? io_r_338_b : _GEN_15317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15319 = 9'h153 == r_count_37_io_out ? io_r_339_b : _GEN_15318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15320 = 9'h154 == r_count_37_io_out ? io_r_340_b : _GEN_15319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15321 = 9'h155 == r_count_37_io_out ? io_r_341_b : _GEN_15320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15322 = 9'h156 == r_count_37_io_out ? io_r_342_b : _GEN_15321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15323 = 9'h157 == r_count_37_io_out ? io_r_343_b : _GEN_15322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15324 = 9'h158 == r_count_37_io_out ? io_r_344_b : _GEN_15323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15325 = 9'h159 == r_count_37_io_out ? io_r_345_b : _GEN_15324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15326 = 9'h15a == r_count_37_io_out ? io_r_346_b : _GEN_15325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15327 = 9'h15b == r_count_37_io_out ? io_r_347_b : _GEN_15326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15328 = 9'h15c == r_count_37_io_out ? io_r_348_b : _GEN_15327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15329 = 9'h15d == r_count_37_io_out ? io_r_349_b : _GEN_15328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15330 = 9'h15e == r_count_37_io_out ? io_r_350_b : _GEN_15329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15331 = 9'h15f == r_count_37_io_out ? io_r_351_b : _GEN_15330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15332 = 9'h160 == r_count_37_io_out ? io_r_352_b : _GEN_15331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15333 = 9'h161 == r_count_37_io_out ? io_r_353_b : _GEN_15332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15334 = 9'h162 == r_count_37_io_out ? io_r_354_b : _GEN_15333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15335 = 9'h163 == r_count_37_io_out ? io_r_355_b : _GEN_15334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15336 = 9'h164 == r_count_37_io_out ? io_r_356_b : _GEN_15335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15337 = 9'h165 == r_count_37_io_out ? io_r_357_b : _GEN_15336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15338 = 9'h166 == r_count_37_io_out ? io_r_358_b : _GEN_15337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15339 = 9'h167 == r_count_37_io_out ? io_r_359_b : _GEN_15338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15340 = 9'h168 == r_count_37_io_out ? io_r_360_b : _GEN_15339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15341 = 9'h169 == r_count_37_io_out ? io_r_361_b : _GEN_15340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15342 = 9'h16a == r_count_37_io_out ? io_r_362_b : _GEN_15341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15343 = 9'h16b == r_count_37_io_out ? io_r_363_b : _GEN_15342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15344 = 9'h16c == r_count_37_io_out ? io_r_364_b : _GEN_15343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15345 = 9'h16d == r_count_37_io_out ? io_r_365_b : _GEN_15344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15346 = 9'h16e == r_count_37_io_out ? io_r_366_b : _GEN_15345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15347 = 9'h16f == r_count_37_io_out ? io_r_367_b : _GEN_15346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15348 = 9'h170 == r_count_37_io_out ? io_r_368_b : _GEN_15347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15349 = 9'h171 == r_count_37_io_out ? io_r_369_b : _GEN_15348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15350 = 9'h172 == r_count_37_io_out ? io_r_370_b : _GEN_15349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15351 = 9'h173 == r_count_37_io_out ? io_r_371_b : _GEN_15350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15352 = 9'h174 == r_count_37_io_out ? io_r_372_b : _GEN_15351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15353 = 9'h175 == r_count_37_io_out ? io_r_373_b : _GEN_15352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15354 = 9'h176 == r_count_37_io_out ? io_r_374_b : _GEN_15353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15355 = 9'h177 == r_count_37_io_out ? io_r_375_b : _GEN_15354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15356 = 9'h178 == r_count_37_io_out ? io_r_376_b : _GEN_15355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15357 = 9'h179 == r_count_37_io_out ? io_r_377_b : _GEN_15356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15358 = 9'h17a == r_count_37_io_out ? io_r_378_b : _GEN_15357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15359 = 9'h17b == r_count_37_io_out ? io_r_379_b : _GEN_15358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15360 = 9'h17c == r_count_37_io_out ? io_r_380_b : _GEN_15359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15361 = 9'h17d == r_count_37_io_out ? io_r_381_b : _GEN_15360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15362 = 9'h17e == r_count_37_io_out ? io_r_382_b : _GEN_15361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15363 = 9'h17f == r_count_37_io_out ? io_r_383_b : _GEN_15362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15364 = 9'h180 == r_count_37_io_out ? io_r_384_b : _GEN_15363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15365 = 9'h181 == r_count_37_io_out ? io_r_385_b : _GEN_15364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15366 = 9'h182 == r_count_37_io_out ? io_r_386_b : _GEN_15365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15367 = 9'h183 == r_count_37_io_out ? io_r_387_b : _GEN_15366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15368 = 9'h184 == r_count_37_io_out ? io_r_388_b : _GEN_15367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15369 = 9'h185 == r_count_37_io_out ? io_r_389_b : _GEN_15368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15370 = 9'h186 == r_count_37_io_out ? io_r_390_b : _GEN_15369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15371 = 9'h187 == r_count_37_io_out ? io_r_391_b : _GEN_15370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15372 = 9'h188 == r_count_37_io_out ? io_r_392_b : _GEN_15371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15373 = 9'h189 == r_count_37_io_out ? io_r_393_b : _GEN_15372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15374 = 9'h18a == r_count_37_io_out ? io_r_394_b : _GEN_15373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15375 = 9'h18b == r_count_37_io_out ? io_r_395_b : _GEN_15374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15376 = 9'h18c == r_count_37_io_out ? io_r_396_b : _GEN_15375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15377 = 9'h18d == r_count_37_io_out ? io_r_397_b : _GEN_15376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15378 = 9'h18e == r_count_37_io_out ? io_r_398_b : _GEN_15377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15381 = 9'h1 == r_count_38_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15382 = 9'h2 == r_count_38_io_out ? io_r_2_b : _GEN_15381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15383 = 9'h3 == r_count_38_io_out ? io_r_3_b : _GEN_15382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15384 = 9'h4 == r_count_38_io_out ? io_r_4_b : _GEN_15383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15385 = 9'h5 == r_count_38_io_out ? io_r_5_b : _GEN_15384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15386 = 9'h6 == r_count_38_io_out ? io_r_6_b : _GEN_15385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15387 = 9'h7 == r_count_38_io_out ? io_r_7_b : _GEN_15386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15388 = 9'h8 == r_count_38_io_out ? io_r_8_b : _GEN_15387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15389 = 9'h9 == r_count_38_io_out ? io_r_9_b : _GEN_15388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15390 = 9'ha == r_count_38_io_out ? io_r_10_b : _GEN_15389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15391 = 9'hb == r_count_38_io_out ? io_r_11_b : _GEN_15390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15392 = 9'hc == r_count_38_io_out ? io_r_12_b : _GEN_15391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15393 = 9'hd == r_count_38_io_out ? io_r_13_b : _GEN_15392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15394 = 9'he == r_count_38_io_out ? io_r_14_b : _GEN_15393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15395 = 9'hf == r_count_38_io_out ? io_r_15_b : _GEN_15394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15396 = 9'h10 == r_count_38_io_out ? io_r_16_b : _GEN_15395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15397 = 9'h11 == r_count_38_io_out ? io_r_17_b : _GEN_15396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15398 = 9'h12 == r_count_38_io_out ? io_r_18_b : _GEN_15397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15399 = 9'h13 == r_count_38_io_out ? io_r_19_b : _GEN_15398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15400 = 9'h14 == r_count_38_io_out ? io_r_20_b : _GEN_15399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15401 = 9'h15 == r_count_38_io_out ? io_r_21_b : _GEN_15400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15402 = 9'h16 == r_count_38_io_out ? io_r_22_b : _GEN_15401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15403 = 9'h17 == r_count_38_io_out ? io_r_23_b : _GEN_15402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15404 = 9'h18 == r_count_38_io_out ? io_r_24_b : _GEN_15403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15405 = 9'h19 == r_count_38_io_out ? io_r_25_b : _GEN_15404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15406 = 9'h1a == r_count_38_io_out ? io_r_26_b : _GEN_15405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15407 = 9'h1b == r_count_38_io_out ? io_r_27_b : _GEN_15406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15408 = 9'h1c == r_count_38_io_out ? io_r_28_b : _GEN_15407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15409 = 9'h1d == r_count_38_io_out ? io_r_29_b : _GEN_15408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15410 = 9'h1e == r_count_38_io_out ? io_r_30_b : _GEN_15409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15411 = 9'h1f == r_count_38_io_out ? io_r_31_b : _GEN_15410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15412 = 9'h20 == r_count_38_io_out ? io_r_32_b : _GEN_15411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15413 = 9'h21 == r_count_38_io_out ? io_r_33_b : _GEN_15412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15414 = 9'h22 == r_count_38_io_out ? io_r_34_b : _GEN_15413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15415 = 9'h23 == r_count_38_io_out ? io_r_35_b : _GEN_15414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15416 = 9'h24 == r_count_38_io_out ? io_r_36_b : _GEN_15415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15417 = 9'h25 == r_count_38_io_out ? io_r_37_b : _GEN_15416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15418 = 9'h26 == r_count_38_io_out ? io_r_38_b : _GEN_15417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15419 = 9'h27 == r_count_38_io_out ? io_r_39_b : _GEN_15418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15420 = 9'h28 == r_count_38_io_out ? io_r_40_b : _GEN_15419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15421 = 9'h29 == r_count_38_io_out ? io_r_41_b : _GEN_15420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15422 = 9'h2a == r_count_38_io_out ? io_r_42_b : _GEN_15421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15423 = 9'h2b == r_count_38_io_out ? io_r_43_b : _GEN_15422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15424 = 9'h2c == r_count_38_io_out ? io_r_44_b : _GEN_15423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15425 = 9'h2d == r_count_38_io_out ? io_r_45_b : _GEN_15424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15426 = 9'h2e == r_count_38_io_out ? io_r_46_b : _GEN_15425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15427 = 9'h2f == r_count_38_io_out ? io_r_47_b : _GEN_15426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15428 = 9'h30 == r_count_38_io_out ? io_r_48_b : _GEN_15427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15429 = 9'h31 == r_count_38_io_out ? io_r_49_b : _GEN_15428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15430 = 9'h32 == r_count_38_io_out ? io_r_50_b : _GEN_15429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15431 = 9'h33 == r_count_38_io_out ? io_r_51_b : _GEN_15430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15432 = 9'h34 == r_count_38_io_out ? io_r_52_b : _GEN_15431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15433 = 9'h35 == r_count_38_io_out ? io_r_53_b : _GEN_15432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15434 = 9'h36 == r_count_38_io_out ? io_r_54_b : _GEN_15433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15435 = 9'h37 == r_count_38_io_out ? io_r_55_b : _GEN_15434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15436 = 9'h38 == r_count_38_io_out ? io_r_56_b : _GEN_15435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15437 = 9'h39 == r_count_38_io_out ? io_r_57_b : _GEN_15436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15438 = 9'h3a == r_count_38_io_out ? io_r_58_b : _GEN_15437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15439 = 9'h3b == r_count_38_io_out ? io_r_59_b : _GEN_15438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15440 = 9'h3c == r_count_38_io_out ? io_r_60_b : _GEN_15439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15441 = 9'h3d == r_count_38_io_out ? io_r_61_b : _GEN_15440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15442 = 9'h3e == r_count_38_io_out ? io_r_62_b : _GEN_15441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15443 = 9'h3f == r_count_38_io_out ? io_r_63_b : _GEN_15442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15444 = 9'h40 == r_count_38_io_out ? io_r_64_b : _GEN_15443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15445 = 9'h41 == r_count_38_io_out ? io_r_65_b : _GEN_15444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15446 = 9'h42 == r_count_38_io_out ? io_r_66_b : _GEN_15445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15447 = 9'h43 == r_count_38_io_out ? io_r_67_b : _GEN_15446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15448 = 9'h44 == r_count_38_io_out ? io_r_68_b : _GEN_15447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15449 = 9'h45 == r_count_38_io_out ? io_r_69_b : _GEN_15448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15450 = 9'h46 == r_count_38_io_out ? io_r_70_b : _GEN_15449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15451 = 9'h47 == r_count_38_io_out ? io_r_71_b : _GEN_15450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15452 = 9'h48 == r_count_38_io_out ? io_r_72_b : _GEN_15451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15453 = 9'h49 == r_count_38_io_out ? io_r_73_b : _GEN_15452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15454 = 9'h4a == r_count_38_io_out ? io_r_74_b : _GEN_15453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15455 = 9'h4b == r_count_38_io_out ? io_r_75_b : _GEN_15454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15456 = 9'h4c == r_count_38_io_out ? io_r_76_b : _GEN_15455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15457 = 9'h4d == r_count_38_io_out ? io_r_77_b : _GEN_15456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15458 = 9'h4e == r_count_38_io_out ? io_r_78_b : _GEN_15457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15459 = 9'h4f == r_count_38_io_out ? io_r_79_b : _GEN_15458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15460 = 9'h50 == r_count_38_io_out ? io_r_80_b : _GEN_15459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15461 = 9'h51 == r_count_38_io_out ? io_r_81_b : _GEN_15460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15462 = 9'h52 == r_count_38_io_out ? io_r_82_b : _GEN_15461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15463 = 9'h53 == r_count_38_io_out ? io_r_83_b : _GEN_15462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15464 = 9'h54 == r_count_38_io_out ? io_r_84_b : _GEN_15463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15465 = 9'h55 == r_count_38_io_out ? io_r_85_b : _GEN_15464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15466 = 9'h56 == r_count_38_io_out ? io_r_86_b : _GEN_15465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15467 = 9'h57 == r_count_38_io_out ? io_r_87_b : _GEN_15466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15468 = 9'h58 == r_count_38_io_out ? io_r_88_b : _GEN_15467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15469 = 9'h59 == r_count_38_io_out ? io_r_89_b : _GEN_15468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15470 = 9'h5a == r_count_38_io_out ? io_r_90_b : _GEN_15469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15471 = 9'h5b == r_count_38_io_out ? io_r_91_b : _GEN_15470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15472 = 9'h5c == r_count_38_io_out ? io_r_92_b : _GEN_15471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15473 = 9'h5d == r_count_38_io_out ? io_r_93_b : _GEN_15472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15474 = 9'h5e == r_count_38_io_out ? io_r_94_b : _GEN_15473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15475 = 9'h5f == r_count_38_io_out ? io_r_95_b : _GEN_15474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15476 = 9'h60 == r_count_38_io_out ? io_r_96_b : _GEN_15475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15477 = 9'h61 == r_count_38_io_out ? io_r_97_b : _GEN_15476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15478 = 9'h62 == r_count_38_io_out ? io_r_98_b : _GEN_15477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15479 = 9'h63 == r_count_38_io_out ? io_r_99_b : _GEN_15478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15480 = 9'h64 == r_count_38_io_out ? io_r_100_b : _GEN_15479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15481 = 9'h65 == r_count_38_io_out ? io_r_101_b : _GEN_15480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15482 = 9'h66 == r_count_38_io_out ? io_r_102_b : _GEN_15481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15483 = 9'h67 == r_count_38_io_out ? io_r_103_b : _GEN_15482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15484 = 9'h68 == r_count_38_io_out ? io_r_104_b : _GEN_15483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15485 = 9'h69 == r_count_38_io_out ? io_r_105_b : _GEN_15484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15486 = 9'h6a == r_count_38_io_out ? io_r_106_b : _GEN_15485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15487 = 9'h6b == r_count_38_io_out ? io_r_107_b : _GEN_15486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15488 = 9'h6c == r_count_38_io_out ? io_r_108_b : _GEN_15487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15489 = 9'h6d == r_count_38_io_out ? io_r_109_b : _GEN_15488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15490 = 9'h6e == r_count_38_io_out ? io_r_110_b : _GEN_15489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15491 = 9'h6f == r_count_38_io_out ? io_r_111_b : _GEN_15490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15492 = 9'h70 == r_count_38_io_out ? io_r_112_b : _GEN_15491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15493 = 9'h71 == r_count_38_io_out ? io_r_113_b : _GEN_15492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15494 = 9'h72 == r_count_38_io_out ? io_r_114_b : _GEN_15493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15495 = 9'h73 == r_count_38_io_out ? io_r_115_b : _GEN_15494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15496 = 9'h74 == r_count_38_io_out ? io_r_116_b : _GEN_15495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15497 = 9'h75 == r_count_38_io_out ? io_r_117_b : _GEN_15496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15498 = 9'h76 == r_count_38_io_out ? io_r_118_b : _GEN_15497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15499 = 9'h77 == r_count_38_io_out ? io_r_119_b : _GEN_15498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15500 = 9'h78 == r_count_38_io_out ? io_r_120_b : _GEN_15499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15501 = 9'h79 == r_count_38_io_out ? io_r_121_b : _GEN_15500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15502 = 9'h7a == r_count_38_io_out ? io_r_122_b : _GEN_15501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15503 = 9'h7b == r_count_38_io_out ? io_r_123_b : _GEN_15502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15504 = 9'h7c == r_count_38_io_out ? io_r_124_b : _GEN_15503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15505 = 9'h7d == r_count_38_io_out ? io_r_125_b : _GEN_15504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15506 = 9'h7e == r_count_38_io_out ? io_r_126_b : _GEN_15505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15507 = 9'h7f == r_count_38_io_out ? io_r_127_b : _GEN_15506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15508 = 9'h80 == r_count_38_io_out ? io_r_128_b : _GEN_15507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15509 = 9'h81 == r_count_38_io_out ? io_r_129_b : _GEN_15508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15510 = 9'h82 == r_count_38_io_out ? io_r_130_b : _GEN_15509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15511 = 9'h83 == r_count_38_io_out ? io_r_131_b : _GEN_15510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15512 = 9'h84 == r_count_38_io_out ? io_r_132_b : _GEN_15511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15513 = 9'h85 == r_count_38_io_out ? io_r_133_b : _GEN_15512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15514 = 9'h86 == r_count_38_io_out ? io_r_134_b : _GEN_15513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15515 = 9'h87 == r_count_38_io_out ? io_r_135_b : _GEN_15514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15516 = 9'h88 == r_count_38_io_out ? io_r_136_b : _GEN_15515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15517 = 9'h89 == r_count_38_io_out ? io_r_137_b : _GEN_15516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15518 = 9'h8a == r_count_38_io_out ? io_r_138_b : _GEN_15517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15519 = 9'h8b == r_count_38_io_out ? io_r_139_b : _GEN_15518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15520 = 9'h8c == r_count_38_io_out ? io_r_140_b : _GEN_15519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15521 = 9'h8d == r_count_38_io_out ? io_r_141_b : _GEN_15520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15522 = 9'h8e == r_count_38_io_out ? io_r_142_b : _GEN_15521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15523 = 9'h8f == r_count_38_io_out ? io_r_143_b : _GEN_15522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15524 = 9'h90 == r_count_38_io_out ? io_r_144_b : _GEN_15523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15525 = 9'h91 == r_count_38_io_out ? io_r_145_b : _GEN_15524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15526 = 9'h92 == r_count_38_io_out ? io_r_146_b : _GEN_15525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15527 = 9'h93 == r_count_38_io_out ? io_r_147_b : _GEN_15526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15528 = 9'h94 == r_count_38_io_out ? io_r_148_b : _GEN_15527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15529 = 9'h95 == r_count_38_io_out ? io_r_149_b : _GEN_15528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15530 = 9'h96 == r_count_38_io_out ? io_r_150_b : _GEN_15529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15531 = 9'h97 == r_count_38_io_out ? io_r_151_b : _GEN_15530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15532 = 9'h98 == r_count_38_io_out ? io_r_152_b : _GEN_15531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15533 = 9'h99 == r_count_38_io_out ? io_r_153_b : _GEN_15532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15534 = 9'h9a == r_count_38_io_out ? io_r_154_b : _GEN_15533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15535 = 9'h9b == r_count_38_io_out ? io_r_155_b : _GEN_15534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15536 = 9'h9c == r_count_38_io_out ? io_r_156_b : _GEN_15535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15537 = 9'h9d == r_count_38_io_out ? io_r_157_b : _GEN_15536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15538 = 9'h9e == r_count_38_io_out ? io_r_158_b : _GEN_15537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15539 = 9'h9f == r_count_38_io_out ? io_r_159_b : _GEN_15538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15540 = 9'ha0 == r_count_38_io_out ? io_r_160_b : _GEN_15539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15541 = 9'ha1 == r_count_38_io_out ? io_r_161_b : _GEN_15540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15542 = 9'ha2 == r_count_38_io_out ? io_r_162_b : _GEN_15541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15543 = 9'ha3 == r_count_38_io_out ? io_r_163_b : _GEN_15542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15544 = 9'ha4 == r_count_38_io_out ? io_r_164_b : _GEN_15543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15545 = 9'ha5 == r_count_38_io_out ? io_r_165_b : _GEN_15544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15546 = 9'ha6 == r_count_38_io_out ? io_r_166_b : _GEN_15545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15547 = 9'ha7 == r_count_38_io_out ? io_r_167_b : _GEN_15546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15548 = 9'ha8 == r_count_38_io_out ? io_r_168_b : _GEN_15547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15549 = 9'ha9 == r_count_38_io_out ? io_r_169_b : _GEN_15548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15550 = 9'haa == r_count_38_io_out ? io_r_170_b : _GEN_15549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15551 = 9'hab == r_count_38_io_out ? io_r_171_b : _GEN_15550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15552 = 9'hac == r_count_38_io_out ? io_r_172_b : _GEN_15551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15553 = 9'had == r_count_38_io_out ? io_r_173_b : _GEN_15552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15554 = 9'hae == r_count_38_io_out ? io_r_174_b : _GEN_15553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15555 = 9'haf == r_count_38_io_out ? io_r_175_b : _GEN_15554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15556 = 9'hb0 == r_count_38_io_out ? io_r_176_b : _GEN_15555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15557 = 9'hb1 == r_count_38_io_out ? io_r_177_b : _GEN_15556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15558 = 9'hb2 == r_count_38_io_out ? io_r_178_b : _GEN_15557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15559 = 9'hb3 == r_count_38_io_out ? io_r_179_b : _GEN_15558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15560 = 9'hb4 == r_count_38_io_out ? io_r_180_b : _GEN_15559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15561 = 9'hb5 == r_count_38_io_out ? io_r_181_b : _GEN_15560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15562 = 9'hb6 == r_count_38_io_out ? io_r_182_b : _GEN_15561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15563 = 9'hb7 == r_count_38_io_out ? io_r_183_b : _GEN_15562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15564 = 9'hb8 == r_count_38_io_out ? io_r_184_b : _GEN_15563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15565 = 9'hb9 == r_count_38_io_out ? io_r_185_b : _GEN_15564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15566 = 9'hba == r_count_38_io_out ? io_r_186_b : _GEN_15565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15567 = 9'hbb == r_count_38_io_out ? io_r_187_b : _GEN_15566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15568 = 9'hbc == r_count_38_io_out ? io_r_188_b : _GEN_15567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15569 = 9'hbd == r_count_38_io_out ? io_r_189_b : _GEN_15568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15570 = 9'hbe == r_count_38_io_out ? io_r_190_b : _GEN_15569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15571 = 9'hbf == r_count_38_io_out ? io_r_191_b : _GEN_15570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15572 = 9'hc0 == r_count_38_io_out ? io_r_192_b : _GEN_15571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15573 = 9'hc1 == r_count_38_io_out ? io_r_193_b : _GEN_15572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15574 = 9'hc2 == r_count_38_io_out ? io_r_194_b : _GEN_15573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15575 = 9'hc3 == r_count_38_io_out ? io_r_195_b : _GEN_15574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15576 = 9'hc4 == r_count_38_io_out ? io_r_196_b : _GEN_15575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15577 = 9'hc5 == r_count_38_io_out ? io_r_197_b : _GEN_15576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15578 = 9'hc6 == r_count_38_io_out ? io_r_198_b : _GEN_15577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15579 = 9'hc7 == r_count_38_io_out ? io_r_199_b : _GEN_15578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15580 = 9'hc8 == r_count_38_io_out ? io_r_200_b : _GEN_15579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15581 = 9'hc9 == r_count_38_io_out ? io_r_201_b : _GEN_15580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15582 = 9'hca == r_count_38_io_out ? io_r_202_b : _GEN_15581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15583 = 9'hcb == r_count_38_io_out ? io_r_203_b : _GEN_15582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15584 = 9'hcc == r_count_38_io_out ? io_r_204_b : _GEN_15583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15585 = 9'hcd == r_count_38_io_out ? io_r_205_b : _GEN_15584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15586 = 9'hce == r_count_38_io_out ? io_r_206_b : _GEN_15585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15587 = 9'hcf == r_count_38_io_out ? io_r_207_b : _GEN_15586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15588 = 9'hd0 == r_count_38_io_out ? io_r_208_b : _GEN_15587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15589 = 9'hd1 == r_count_38_io_out ? io_r_209_b : _GEN_15588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15590 = 9'hd2 == r_count_38_io_out ? io_r_210_b : _GEN_15589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15591 = 9'hd3 == r_count_38_io_out ? io_r_211_b : _GEN_15590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15592 = 9'hd4 == r_count_38_io_out ? io_r_212_b : _GEN_15591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15593 = 9'hd5 == r_count_38_io_out ? io_r_213_b : _GEN_15592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15594 = 9'hd6 == r_count_38_io_out ? io_r_214_b : _GEN_15593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15595 = 9'hd7 == r_count_38_io_out ? io_r_215_b : _GEN_15594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15596 = 9'hd8 == r_count_38_io_out ? io_r_216_b : _GEN_15595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15597 = 9'hd9 == r_count_38_io_out ? io_r_217_b : _GEN_15596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15598 = 9'hda == r_count_38_io_out ? io_r_218_b : _GEN_15597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15599 = 9'hdb == r_count_38_io_out ? io_r_219_b : _GEN_15598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15600 = 9'hdc == r_count_38_io_out ? io_r_220_b : _GEN_15599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15601 = 9'hdd == r_count_38_io_out ? io_r_221_b : _GEN_15600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15602 = 9'hde == r_count_38_io_out ? io_r_222_b : _GEN_15601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15603 = 9'hdf == r_count_38_io_out ? io_r_223_b : _GEN_15602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15604 = 9'he0 == r_count_38_io_out ? io_r_224_b : _GEN_15603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15605 = 9'he1 == r_count_38_io_out ? io_r_225_b : _GEN_15604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15606 = 9'he2 == r_count_38_io_out ? io_r_226_b : _GEN_15605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15607 = 9'he3 == r_count_38_io_out ? io_r_227_b : _GEN_15606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15608 = 9'he4 == r_count_38_io_out ? io_r_228_b : _GEN_15607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15609 = 9'he5 == r_count_38_io_out ? io_r_229_b : _GEN_15608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15610 = 9'he6 == r_count_38_io_out ? io_r_230_b : _GEN_15609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15611 = 9'he7 == r_count_38_io_out ? io_r_231_b : _GEN_15610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15612 = 9'he8 == r_count_38_io_out ? io_r_232_b : _GEN_15611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15613 = 9'he9 == r_count_38_io_out ? io_r_233_b : _GEN_15612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15614 = 9'hea == r_count_38_io_out ? io_r_234_b : _GEN_15613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15615 = 9'heb == r_count_38_io_out ? io_r_235_b : _GEN_15614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15616 = 9'hec == r_count_38_io_out ? io_r_236_b : _GEN_15615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15617 = 9'hed == r_count_38_io_out ? io_r_237_b : _GEN_15616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15618 = 9'hee == r_count_38_io_out ? io_r_238_b : _GEN_15617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15619 = 9'hef == r_count_38_io_out ? io_r_239_b : _GEN_15618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15620 = 9'hf0 == r_count_38_io_out ? io_r_240_b : _GEN_15619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15621 = 9'hf1 == r_count_38_io_out ? io_r_241_b : _GEN_15620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15622 = 9'hf2 == r_count_38_io_out ? io_r_242_b : _GEN_15621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15623 = 9'hf3 == r_count_38_io_out ? io_r_243_b : _GEN_15622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15624 = 9'hf4 == r_count_38_io_out ? io_r_244_b : _GEN_15623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15625 = 9'hf5 == r_count_38_io_out ? io_r_245_b : _GEN_15624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15626 = 9'hf6 == r_count_38_io_out ? io_r_246_b : _GEN_15625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15627 = 9'hf7 == r_count_38_io_out ? io_r_247_b : _GEN_15626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15628 = 9'hf8 == r_count_38_io_out ? io_r_248_b : _GEN_15627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15629 = 9'hf9 == r_count_38_io_out ? io_r_249_b : _GEN_15628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15630 = 9'hfa == r_count_38_io_out ? io_r_250_b : _GEN_15629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15631 = 9'hfb == r_count_38_io_out ? io_r_251_b : _GEN_15630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15632 = 9'hfc == r_count_38_io_out ? io_r_252_b : _GEN_15631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15633 = 9'hfd == r_count_38_io_out ? io_r_253_b : _GEN_15632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15634 = 9'hfe == r_count_38_io_out ? io_r_254_b : _GEN_15633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15635 = 9'hff == r_count_38_io_out ? io_r_255_b : _GEN_15634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15636 = 9'h100 == r_count_38_io_out ? io_r_256_b : _GEN_15635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15637 = 9'h101 == r_count_38_io_out ? io_r_257_b : _GEN_15636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15638 = 9'h102 == r_count_38_io_out ? io_r_258_b : _GEN_15637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15639 = 9'h103 == r_count_38_io_out ? io_r_259_b : _GEN_15638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15640 = 9'h104 == r_count_38_io_out ? io_r_260_b : _GEN_15639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15641 = 9'h105 == r_count_38_io_out ? io_r_261_b : _GEN_15640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15642 = 9'h106 == r_count_38_io_out ? io_r_262_b : _GEN_15641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15643 = 9'h107 == r_count_38_io_out ? io_r_263_b : _GEN_15642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15644 = 9'h108 == r_count_38_io_out ? io_r_264_b : _GEN_15643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15645 = 9'h109 == r_count_38_io_out ? io_r_265_b : _GEN_15644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15646 = 9'h10a == r_count_38_io_out ? io_r_266_b : _GEN_15645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15647 = 9'h10b == r_count_38_io_out ? io_r_267_b : _GEN_15646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15648 = 9'h10c == r_count_38_io_out ? io_r_268_b : _GEN_15647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15649 = 9'h10d == r_count_38_io_out ? io_r_269_b : _GEN_15648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15650 = 9'h10e == r_count_38_io_out ? io_r_270_b : _GEN_15649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15651 = 9'h10f == r_count_38_io_out ? io_r_271_b : _GEN_15650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15652 = 9'h110 == r_count_38_io_out ? io_r_272_b : _GEN_15651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15653 = 9'h111 == r_count_38_io_out ? io_r_273_b : _GEN_15652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15654 = 9'h112 == r_count_38_io_out ? io_r_274_b : _GEN_15653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15655 = 9'h113 == r_count_38_io_out ? io_r_275_b : _GEN_15654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15656 = 9'h114 == r_count_38_io_out ? io_r_276_b : _GEN_15655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15657 = 9'h115 == r_count_38_io_out ? io_r_277_b : _GEN_15656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15658 = 9'h116 == r_count_38_io_out ? io_r_278_b : _GEN_15657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15659 = 9'h117 == r_count_38_io_out ? io_r_279_b : _GEN_15658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15660 = 9'h118 == r_count_38_io_out ? io_r_280_b : _GEN_15659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15661 = 9'h119 == r_count_38_io_out ? io_r_281_b : _GEN_15660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15662 = 9'h11a == r_count_38_io_out ? io_r_282_b : _GEN_15661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15663 = 9'h11b == r_count_38_io_out ? io_r_283_b : _GEN_15662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15664 = 9'h11c == r_count_38_io_out ? io_r_284_b : _GEN_15663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15665 = 9'h11d == r_count_38_io_out ? io_r_285_b : _GEN_15664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15666 = 9'h11e == r_count_38_io_out ? io_r_286_b : _GEN_15665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15667 = 9'h11f == r_count_38_io_out ? io_r_287_b : _GEN_15666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15668 = 9'h120 == r_count_38_io_out ? io_r_288_b : _GEN_15667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15669 = 9'h121 == r_count_38_io_out ? io_r_289_b : _GEN_15668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15670 = 9'h122 == r_count_38_io_out ? io_r_290_b : _GEN_15669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15671 = 9'h123 == r_count_38_io_out ? io_r_291_b : _GEN_15670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15672 = 9'h124 == r_count_38_io_out ? io_r_292_b : _GEN_15671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15673 = 9'h125 == r_count_38_io_out ? io_r_293_b : _GEN_15672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15674 = 9'h126 == r_count_38_io_out ? io_r_294_b : _GEN_15673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15675 = 9'h127 == r_count_38_io_out ? io_r_295_b : _GEN_15674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15676 = 9'h128 == r_count_38_io_out ? io_r_296_b : _GEN_15675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15677 = 9'h129 == r_count_38_io_out ? io_r_297_b : _GEN_15676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15678 = 9'h12a == r_count_38_io_out ? io_r_298_b : _GEN_15677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15679 = 9'h12b == r_count_38_io_out ? io_r_299_b : _GEN_15678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15680 = 9'h12c == r_count_38_io_out ? io_r_300_b : _GEN_15679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15681 = 9'h12d == r_count_38_io_out ? io_r_301_b : _GEN_15680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15682 = 9'h12e == r_count_38_io_out ? io_r_302_b : _GEN_15681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15683 = 9'h12f == r_count_38_io_out ? io_r_303_b : _GEN_15682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15684 = 9'h130 == r_count_38_io_out ? io_r_304_b : _GEN_15683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15685 = 9'h131 == r_count_38_io_out ? io_r_305_b : _GEN_15684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15686 = 9'h132 == r_count_38_io_out ? io_r_306_b : _GEN_15685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15687 = 9'h133 == r_count_38_io_out ? io_r_307_b : _GEN_15686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15688 = 9'h134 == r_count_38_io_out ? io_r_308_b : _GEN_15687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15689 = 9'h135 == r_count_38_io_out ? io_r_309_b : _GEN_15688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15690 = 9'h136 == r_count_38_io_out ? io_r_310_b : _GEN_15689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15691 = 9'h137 == r_count_38_io_out ? io_r_311_b : _GEN_15690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15692 = 9'h138 == r_count_38_io_out ? io_r_312_b : _GEN_15691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15693 = 9'h139 == r_count_38_io_out ? io_r_313_b : _GEN_15692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15694 = 9'h13a == r_count_38_io_out ? io_r_314_b : _GEN_15693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15695 = 9'h13b == r_count_38_io_out ? io_r_315_b : _GEN_15694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15696 = 9'h13c == r_count_38_io_out ? io_r_316_b : _GEN_15695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15697 = 9'h13d == r_count_38_io_out ? io_r_317_b : _GEN_15696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15698 = 9'h13e == r_count_38_io_out ? io_r_318_b : _GEN_15697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15699 = 9'h13f == r_count_38_io_out ? io_r_319_b : _GEN_15698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15700 = 9'h140 == r_count_38_io_out ? io_r_320_b : _GEN_15699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15701 = 9'h141 == r_count_38_io_out ? io_r_321_b : _GEN_15700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15702 = 9'h142 == r_count_38_io_out ? io_r_322_b : _GEN_15701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15703 = 9'h143 == r_count_38_io_out ? io_r_323_b : _GEN_15702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15704 = 9'h144 == r_count_38_io_out ? io_r_324_b : _GEN_15703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15705 = 9'h145 == r_count_38_io_out ? io_r_325_b : _GEN_15704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15706 = 9'h146 == r_count_38_io_out ? io_r_326_b : _GEN_15705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15707 = 9'h147 == r_count_38_io_out ? io_r_327_b : _GEN_15706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15708 = 9'h148 == r_count_38_io_out ? io_r_328_b : _GEN_15707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15709 = 9'h149 == r_count_38_io_out ? io_r_329_b : _GEN_15708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15710 = 9'h14a == r_count_38_io_out ? io_r_330_b : _GEN_15709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15711 = 9'h14b == r_count_38_io_out ? io_r_331_b : _GEN_15710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15712 = 9'h14c == r_count_38_io_out ? io_r_332_b : _GEN_15711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15713 = 9'h14d == r_count_38_io_out ? io_r_333_b : _GEN_15712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15714 = 9'h14e == r_count_38_io_out ? io_r_334_b : _GEN_15713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15715 = 9'h14f == r_count_38_io_out ? io_r_335_b : _GEN_15714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15716 = 9'h150 == r_count_38_io_out ? io_r_336_b : _GEN_15715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15717 = 9'h151 == r_count_38_io_out ? io_r_337_b : _GEN_15716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15718 = 9'h152 == r_count_38_io_out ? io_r_338_b : _GEN_15717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15719 = 9'h153 == r_count_38_io_out ? io_r_339_b : _GEN_15718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15720 = 9'h154 == r_count_38_io_out ? io_r_340_b : _GEN_15719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15721 = 9'h155 == r_count_38_io_out ? io_r_341_b : _GEN_15720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15722 = 9'h156 == r_count_38_io_out ? io_r_342_b : _GEN_15721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15723 = 9'h157 == r_count_38_io_out ? io_r_343_b : _GEN_15722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15724 = 9'h158 == r_count_38_io_out ? io_r_344_b : _GEN_15723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15725 = 9'h159 == r_count_38_io_out ? io_r_345_b : _GEN_15724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15726 = 9'h15a == r_count_38_io_out ? io_r_346_b : _GEN_15725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15727 = 9'h15b == r_count_38_io_out ? io_r_347_b : _GEN_15726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15728 = 9'h15c == r_count_38_io_out ? io_r_348_b : _GEN_15727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15729 = 9'h15d == r_count_38_io_out ? io_r_349_b : _GEN_15728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15730 = 9'h15e == r_count_38_io_out ? io_r_350_b : _GEN_15729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15731 = 9'h15f == r_count_38_io_out ? io_r_351_b : _GEN_15730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15732 = 9'h160 == r_count_38_io_out ? io_r_352_b : _GEN_15731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15733 = 9'h161 == r_count_38_io_out ? io_r_353_b : _GEN_15732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15734 = 9'h162 == r_count_38_io_out ? io_r_354_b : _GEN_15733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15735 = 9'h163 == r_count_38_io_out ? io_r_355_b : _GEN_15734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15736 = 9'h164 == r_count_38_io_out ? io_r_356_b : _GEN_15735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15737 = 9'h165 == r_count_38_io_out ? io_r_357_b : _GEN_15736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15738 = 9'h166 == r_count_38_io_out ? io_r_358_b : _GEN_15737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15739 = 9'h167 == r_count_38_io_out ? io_r_359_b : _GEN_15738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15740 = 9'h168 == r_count_38_io_out ? io_r_360_b : _GEN_15739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15741 = 9'h169 == r_count_38_io_out ? io_r_361_b : _GEN_15740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15742 = 9'h16a == r_count_38_io_out ? io_r_362_b : _GEN_15741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15743 = 9'h16b == r_count_38_io_out ? io_r_363_b : _GEN_15742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15744 = 9'h16c == r_count_38_io_out ? io_r_364_b : _GEN_15743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15745 = 9'h16d == r_count_38_io_out ? io_r_365_b : _GEN_15744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15746 = 9'h16e == r_count_38_io_out ? io_r_366_b : _GEN_15745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15747 = 9'h16f == r_count_38_io_out ? io_r_367_b : _GEN_15746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15748 = 9'h170 == r_count_38_io_out ? io_r_368_b : _GEN_15747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15749 = 9'h171 == r_count_38_io_out ? io_r_369_b : _GEN_15748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15750 = 9'h172 == r_count_38_io_out ? io_r_370_b : _GEN_15749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15751 = 9'h173 == r_count_38_io_out ? io_r_371_b : _GEN_15750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15752 = 9'h174 == r_count_38_io_out ? io_r_372_b : _GEN_15751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15753 = 9'h175 == r_count_38_io_out ? io_r_373_b : _GEN_15752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15754 = 9'h176 == r_count_38_io_out ? io_r_374_b : _GEN_15753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15755 = 9'h177 == r_count_38_io_out ? io_r_375_b : _GEN_15754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15756 = 9'h178 == r_count_38_io_out ? io_r_376_b : _GEN_15755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15757 = 9'h179 == r_count_38_io_out ? io_r_377_b : _GEN_15756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15758 = 9'h17a == r_count_38_io_out ? io_r_378_b : _GEN_15757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15759 = 9'h17b == r_count_38_io_out ? io_r_379_b : _GEN_15758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15760 = 9'h17c == r_count_38_io_out ? io_r_380_b : _GEN_15759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15761 = 9'h17d == r_count_38_io_out ? io_r_381_b : _GEN_15760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15762 = 9'h17e == r_count_38_io_out ? io_r_382_b : _GEN_15761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15763 = 9'h17f == r_count_38_io_out ? io_r_383_b : _GEN_15762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15764 = 9'h180 == r_count_38_io_out ? io_r_384_b : _GEN_15763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15765 = 9'h181 == r_count_38_io_out ? io_r_385_b : _GEN_15764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15766 = 9'h182 == r_count_38_io_out ? io_r_386_b : _GEN_15765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15767 = 9'h183 == r_count_38_io_out ? io_r_387_b : _GEN_15766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15768 = 9'h184 == r_count_38_io_out ? io_r_388_b : _GEN_15767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15769 = 9'h185 == r_count_38_io_out ? io_r_389_b : _GEN_15768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15770 = 9'h186 == r_count_38_io_out ? io_r_390_b : _GEN_15769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15771 = 9'h187 == r_count_38_io_out ? io_r_391_b : _GEN_15770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15772 = 9'h188 == r_count_38_io_out ? io_r_392_b : _GEN_15771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15773 = 9'h189 == r_count_38_io_out ? io_r_393_b : _GEN_15772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15774 = 9'h18a == r_count_38_io_out ? io_r_394_b : _GEN_15773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15775 = 9'h18b == r_count_38_io_out ? io_r_395_b : _GEN_15774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15776 = 9'h18c == r_count_38_io_out ? io_r_396_b : _GEN_15775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15777 = 9'h18d == r_count_38_io_out ? io_r_397_b : _GEN_15776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15778 = 9'h18e == r_count_38_io_out ? io_r_398_b : _GEN_15777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15781 = 9'h1 == r_count_39_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15782 = 9'h2 == r_count_39_io_out ? io_r_2_b : _GEN_15781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15783 = 9'h3 == r_count_39_io_out ? io_r_3_b : _GEN_15782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15784 = 9'h4 == r_count_39_io_out ? io_r_4_b : _GEN_15783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15785 = 9'h5 == r_count_39_io_out ? io_r_5_b : _GEN_15784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15786 = 9'h6 == r_count_39_io_out ? io_r_6_b : _GEN_15785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15787 = 9'h7 == r_count_39_io_out ? io_r_7_b : _GEN_15786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15788 = 9'h8 == r_count_39_io_out ? io_r_8_b : _GEN_15787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15789 = 9'h9 == r_count_39_io_out ? io_r_9_b : _GEN_15788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15790 = 9'ha == r_count_39_io_out ? io_r_10_b : _GEN_15789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15791 = 9'hb == r_count_39_io_out ? io_r_11_b : _GEN_15790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15792 = 9'hc == r_count_39_io_out ? io_r_12_b : _GEN_15791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15793 = 9'hd == r_count_39_io_out ? io_r_13_b : _GEN_15792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15794 = 9'he == r_count_39_io_out ? io_r_14_b : _GEN_15793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15795 = 9'hf == r_count_39_io_out ? io_r_15_b : _GEN_15794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15796 = 9'h10 == r_count_39_io_out ? io_r_16_b : _GEN_15795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15797 = 9'h11 == r_count_39_io_out ? io_r_17_b : _GEN_15796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15798 = 9'h12 == r_count_39_io_out ? io_r_18_b : _GEN_15797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15799 = 9'h13 == r_count_39_io_out ? io_r_19_b : _GEN_15798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15800 = 9'h14 == r_count_39_io_out ? io_r_20_b : _GEN_15799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15801 = 9'h15 == r_count_39_io_out ? io_r_21_b : _GEN_15800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15802 = 9'h16 == r_count_39_io_out ? io_r_22_b : _GEN_15801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15803 = 9'h17 == r_count_39_io_out ? io_r_23_b : _GEN_15802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15804 = 9'h18 == r_count_39_io_out ? io_r_24_b : _GEN_15803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15805 = 9'h19 == r_count_39_io_out ? io_r_25_b : _GEN_15804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15806 = 9'h1a == r_count_39_io_out ? io_r_26_b : _GEN_15805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15807 = 9'h1b == r_count_39_io_out ? io_r_27_b : _GEN_15806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15808 = 9'h1c == r_count_39_io_out ? io_r_28_b : _GEN_15807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15809 = 9'h1d == r_count_39_io_out ? io_r_29_b : _GEN_15808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15810 = 9'h1e == r_count_39_io_out ? io_r_30_b : _GEN_15809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15811 = 9'h1f == r_count_39_io_out ? io_r_31_b : _GEN_15810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15812 = 9'h20 == r_count_39_io_out ? io_r_32_b : _GEN_15811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15813 = 9'h21 == r_count_39_io_out ? io_r_33_b : _GEN_15812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15814 = 9'h22 == r_count_39_io_out ? io_r_34_b : _GEN_15813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15815 = 9'h23 == r_count_39_io_out ? io_r_35_b : _GEN_15814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15816 = 9'h24 == r_count_39_io_out ? io_r_36_b : _GEN_15815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15817 = 9'h25 == r_count_39_io_out ? io_r_37_b : _GEN_15816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15818 = 9'h26 == r_count_39_io_out ? io_r_38_b : _GEN_15817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15819 = 9'h27 == r_count_39_io_out ? io_r_39_b : _GEN_15818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15820 = 9'h28 == r_count_39_io_out ? io_r_40_b : _GEN_15819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15821 = 9'h29 == r_count_39_io_out ? io_r_41_b : _GEN_15820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15822 = 9'h2a == r_count_39_io_out ? io_r_42_b : _GEN_15821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15823 = 9'h2b == r_count_39_io_out ? io_r_43_b : _GEN_15822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15824 = 9'h2c == r_count_39_io_out ? io_r_44_b : _GEN_15823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15825 = 9'h2d == r_count_39_io_out ? io_r_45_b : _GEN_15824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15826 = 9'h2e == r_count_39_io_out ? io_r_46_b : _GEN_15825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15827 = 9'h2f == r_count_39_io_out ? io_r_47_b : _GEN_15826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15828 = 9'h30 == r_count_39_io_out ? io_r_48_b : _GEN_15827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15829 = 9'h31 == r_count_39_io_out ? io_r_49_b : _GEN_15828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15830 = 9'h32 == r_count_39_io_out ? io_r_50_b : _GEN_15829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15831 = 9'h33 == r_count_39_io_out ? io_r_51_b : _GEN_15830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15832 = 9'h34 == r_count_39_io_out ? io_r_52_b : _GEN_15831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15833 = 9'h35 == r_count_39_io_out ? io_r_53_b : _GEN_15832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15834 = 9'h36 == r_count_39_io_out ? io_r_54_b : _GEN_15833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15835 = 9'h37 == r_count_39_io_out ? io_r_55_b : _GEN_15834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15836 = 9'h38 == r_count_39_io_out ? io_r_56_b : _GEN_15835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15837 = 9'h39 == r_count_39_io_out ? io_r_57_b : _GEN_15836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15838 = 9'h3a == r_count_39_io_out ? io_r_58_b : _GEN_15837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15839 = 9'h3b == r_count_39_io_out ? io_r_59_b : _GEN_15838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15840 = 9'h3c == r_count_39_io_out ? io_r_60_b : _GEN_15839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15841 = 9'h3d == r_count_39_io_out ? io_r_61_b : _GEN_15840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15842 = 9'h3e == r_count_39_io_out ? io_r_62_b : _GEN_15841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15843 = 9'h3f == r_count_39_io_out ? io_r_63_b : _GEN_15842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15844 = 9'h40 == r_count_39_io_out ? io_r_64_b : _GEN_15843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15845 = 9'h41 == r_count_39_io_out ? io_r_65_b : _GEN_15844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15846 = 9'h42 == r_count_39_io_out ? io_r_66_b : _GEN_15845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15847 = 9'h43 == r_count_39_io_out ? io_r_67_b : _GEN_15846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15848 = 9'h44 == r_count_39_io_out ? io_r_68_b : _GEN_15847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15849 = 9'h45 == r_count_39_io_out ? io_r_69_b : _GEN_15848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15850 = 9'h46 == r_count_39_io_out ? io_r_70_b : _GEN_15849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15851 = 9'h47 == r_count_39_io_out ? io_r_71_b : _GEN_15850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15852 = 9'h48 == r_count_39_io_out ? io_r_72_b : _GEN_15851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15853 = 9'h49 == r_count_39_io_out ? io_r_73_b : _GEN_15852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15854 = 9'h4a == r_count_39_io_out ? io_r_74_b : _GEN_15853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15855 = 9'h4b == r_count_39_io_out ? io_r_75_b : _GEN_15854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15856 = 9'h4c == r_count_39_io_out ? io_r_76_b : _GEN_15855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15857 = 9'h4d == r_count_39_io_out ? io_r_77_b : _GEN_15856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15858 = 9'h4e == r_count_39_io_out ? io_r_78_b : _GEN_15857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15859 = 9'h4f == r_count_39_io_out ? io_r_79_b : _GEN_15858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15860 = 9'h50 == r_count_39_io_out ? io_r_80_b : _GEN_15859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15861 = 9'h51 == r_count_39_io_out ? io_r_81_b : _GEN_15860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15862 = 9'h52 == r_count_39_io_out ? io_r_82_b : _GEN_15861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15863 = 9'h53 == r_count_39_io_out ? io_r_83_b : _GEN_15862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15864 = 9'h54 == r_count_39_io_out ? io_r_84_b : _GEN_15863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15865 = 9'h55 == r_count_39_io_out ? io_r_85_b : _GEN_15864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15866 = 9'h56 == r_count_39_io_out ? io_r_86_b : _GEN_15865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15867 = 9'h57 == r_count_39_io_out ? io_r_87_b : _GEN_15866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15868 = 9'h58 == r_count_39_io_out ? io_r_88_b : _GEN_15867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15869 = 9'h59 == r_count_39_io_out ? io_r_89_b : _GEN_15868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15870 = 9'h5a == r_count_39_io_out ? io_r_90_b : _GEN_15869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15871 = 9'h5b == r_count_39_io_out ? io_r_91_b : _GEN_15870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15872 = 9'h5c == r_count_39_io_out ? io_r_92_b : _GEN_15871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15873 = 9'h5d == r_count_39_io_out ? io_r_93_b : _GEN_15872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15874 = 9'h5e == r_count_39_io_out ? io_r_94_b : _GEN_15873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15875 = 9'h5f == r_count_39_io_out ? io_r_95_b : _GEN_15874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15876 = 9'h60 == r_count_39_io_out ? io_r_96_b : _GEN_15875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15877 = 9'h61 == r_count_39_io_out ? io_r_97_b : _GEN_15876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15878 = 9'h62 == r_count_39_io_out ? io_r_98_b : _GEN_15877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15879 = 9'h63 == r_count_39_io_out ? io_r_99_b : _GEN_15878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15880 = 9'h64 == r_count_39_io_out ? io_r_100_b : _GEN_15879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15881 = 9'h65 == r_count_39_io_out ? io_r_101_b : _GEN_15880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15882 = 9'h66 == r_count_39_io_out ? io_r_102_b : _GEN_15881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15883 = 9'h67 == r_count_39_io_out ? io_r_103_b : _GEN_15882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15884 = 9'h68 == r_count_39_io_out ? io_r_104_b : _GEN_15883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15885 = 9'h69 == r_count_39_io_out ? io_r_105_b : _GEN_15884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15886 = 9'h6a == r_count_39_io_out ? io_r_106_b : _GEN_15885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15887 = 9'h6b == r_count_39_io_out ? io_r_107_b : _GEN_15886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15888 = 9'h6c == r_count_39_io_out ? io_r_108_b : _GEN_15887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15889 = 9'h6d == r_count_39_io_out ? io_r_109_b : _GEN_15888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15890 = 9'h6e == r_count_39_io_out ? io_r_110_b : _GEN_15889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15891 = 9'h6f == r_count_39_io_out ? io_r_111_b : _GEN_15890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15892 = 9'h70 == r_count_39_io_out ? io_r_112_b : _GEN_15891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15893 = 9'h71 == r_count_39_io_out ? io_r_113_b : _GEN_15892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15894 = 9'h72 == r_count_39_io_out ? io_r_114_b : _GEN_15893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15895 = 9'h73 == r_count_39_io_out ? io_r_115_b : _GEN_15894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15896 = 9'h74 == r_count_39_io_out ? io_r_116_b : _GEN_15895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15897 = 9'h75 == r_count_39_io_out ? io_r_117_b : _GEN_15896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15898 = 9'h76 == r_count_39_io_out ? io_r_118_b : _GEN_15897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15899 = 9'h77 == r_count_39_io_out ? io_r_119_b : _GEN_15898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15900 = 9'h78 == r_count_39_io_out ? io_r_120_b : _GEN_15899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15901 = 9'h79 == r_count_39_io_out ? io_r_121_b : _GEN_15900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15902 = 9'h7a == r_count_39_io_out ? io_r_122_b : _GEN_15901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15903 = 9'h7b == r_count_39_io_out ? io_r_123_b : _GEN_15902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15904 = 9'h7c == r_count_39_io_out ? io_r_124_b : _GEN_15903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15905 = 9'h7d == r_count_39_io_out ? io_r_125_b : _GEN_15904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15906 = 9'h7e == r_count_39_io_out ? io_r_126_b : _GEN_15905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15907 = 9'h7f == r_count_39_io_out ? io_r_127_b : _GEN_15906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15908 = 9'h80 == r_count_39_io_out ? io_r_128_b : _GEN_15907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15909 = 9'h81 == r_count_39_io_out ? io_r_129_b : _GEN_15908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15910 = 9'h82 == r_count_39_io_out ? io_r_130_b : _GEN_15909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15911 = 9'h83 == r_count_39_io_out ? io_r_131_b : _GEN_15910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15912 = 9'h84 == r_count_39_io_out ? io_r_132_b : _GEN_15911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15913 = 9'h85 == r_count_39_io_out ? io_r_133_b : _GEN_15912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15914 = 9'h86 == r_count_39_io_out ? io_r_134_b : _GEN_15913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15915 = 9'h87 == r_count_39_io_out ? io_r_135_b : _GEN_15914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15916 = 9'h88 == r_count_39_io_out ? io_r_136_b : _GEN_15915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15917 = 9'h89 == r_count_39_io_out ? io_r_137_b : _GEN_15916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15918 = 9'h8a == r_count_39_io_out ? io_r_138_b : _GEN_15917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15919 = 9'h8b == r_count_39_io_out ? io_r_139_b : _GEN_15918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15920 = 9'h8c == r_count_39_io_out ? io_r_140_b : _GEN_15919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15921 = 9'h8d == r_count_39_io_out ? io_r_141_b : _GEN_15920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15922 = 9'h8e == r_count_39_io_out ? io_r_142_b : _GEN_15921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15923 = 9'h8f == r_count_39_io_out ? io_r_143_b : _GEN_15922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15924 = 9'h90 == r_count_39_io_out ? io_r_144_b : _GEN_15923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15925 = 9'h91 == r_count_39_io_out ? io_r_145_b : _GEN_15924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15926 = 9'h92 == r_count_39_io_out ? io_r_146_b : _GEN_15925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15927 = 9'h93 == r_count_39_io_out ? io_r_147_b : _GEN_15926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15928 = 9'h94 == r_count_39_io_out ? io_r_148_b : _GEN_15927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15929 = 9'h95 == r_count_39_io_out ? io_r_149_b : _GEN_15928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15930 = 9'h96 == r_count_39_io_out ? io_r_150_b : _GEN_15929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15931 = 9'h97 == r_count_39_io_out ? io_r_151_b : _GEN_15930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15932 = 9'h98 == r_count_39_io_out ? io_r_152_b : _GEN_15931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15933 = 9'h99 == r_count_39_io_out ? io_r_153_b : _GEN_15932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15934 = 9'h9a == r_count_39_io_out ? io_r_154_b : _GEN_15933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15935 = 9'h9b == r_count_39_io_out ? io_r_155_b : _GEN_15934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15936 = 9'h9c == r_count_39_io_out ? io_r_156_b : _GEN_15935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15937 = 9'h9d == r_count_39_io_out ? io_r_157_b : _GEN_15936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15938 = 9'h9e == r_count_39_io_out ? io_r_158_b : _GEN_15937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15939 = 9'h9f == r_count_39_io_out ? io_r_159_b : _GEN_15938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15940 = 9'ha0 == r_count_39_io_out ? io_r_160_b : _GEN_15939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15941 = 9'ha1 == r_count_39_io_out ? io_r_161_b : _GEN_15940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15942 = 9'ha2 == r_count_39_io_out ? io_r_162_b : _GEN_15941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15943 = 9'ha3 == r_count_39_io_out ? io_r_163_b : _GEN_15942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15944 = 9'ha4 == r_count_39_io_out ? io_r_164_b : _GEN_15943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15945 = 9'ha5 == r_count_39_io_out ? io_r_165_b : _GEN_15944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15946 = 9'ha6 == r_count_39_io_out ? io_r_166_b : _GEN_15945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15947 = 9'ha7 == r_count_39_io_out ? io_r_167_b : _GEN_15946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15948 = 9'ha8 == r_count_39_io_out ? io_r_168_b : _GEN_15947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15949 = 9'ha9 == r_count_39_io_out ? io_r_169_b : _GEN_15948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15950 = 9'haa == r_count_39_io_out ? io_r_170_b : _GEN_15949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15951 = 9'hab == r_count_39_io_out ? io_r_171_b : _GEN_15950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15952 = 9'hac == r_count_39_io_out ? io_r_172_b : _GEN_15951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15953 = 9'had == r_count_39_io_out ? io_r_173_b : _GEN_15952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15954 = 9'hae == r_count_39_io_out ? io_r_174_b : _GEN_15953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15955 = 9'haf == r_count_39_io_out ? io_r_175_b : _GEN_15954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15956 = 9'hb0 == r_count_39_io_out ? io_r_176_b : _GEN_15955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15957 = 9'hb1 == r_count_39_io_out ? io_r_177_b : _GEN_15956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15958 = 9'hb2 == r_count_39_io_out ? io_r_178_b : _GEN_15957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15959 = 9'hb3 == r_count_39_io_out ? io_r_179_b : _GEN_15958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15960 = 9'hb4 == r_count_39_io_out ? io_r_180_b : _GEN_15959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15961 = 9'hb5 == r_count_39_io_out ? io_r_181_b : _GEN_15960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15962 = 9'hb6 == r_count_39_io_out ? io_r_182_b : _GEN_15961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15963 = 9'hb7 == r_count_39_io_out ? io_r_183_b : _GEN_15962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15964 = 9'hb8 == r_count_39_io_out ? io_r_184_b : _GEN_15963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15965 = 9'hb9 == r_count_39_io_out ? io_r_185_b : _GEN_15964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15966 = 9'hba == r_count_39_io_out ? io_r_186_b : _GEN_15965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15967 = 9'hbb == r_count_39_io_out ? io_r_187_b : _GEN_15966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15968 = 9'hbc == r_count_39_io_out ? io_r_188_b : _GEN_15967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15969 = 9'hbd == r_count_39_io_out ? io_r_189_b : _GEN_15968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15970 = 9'hbe == r_count_39_io_out ? io_r_190_b : _GEN_15969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15971 = 9'hbf == r_count_39_io_out ? io_r_191_b : _GEN_15970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15972 = 9'hc0 == r_count_39_io_out ? io_r_192_b : _GEN_15971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15973 = 9'hc1 == r_count_39_io_out ? io_r_193_b : _GEN_15972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15974 = 9'hc2 == r_count_39_io_out ? io_r_194_b : _GEN_15973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15975 = 9'hc3 == r_count_39_io_out ? io_r_195_b : _GEN_15974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15976 = 9'hc4 == r_count_39_io_out ? io_r_196_b : _GEN_15975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15977 = 9'hc5 == r_count_39_io_out ? io_r_197_b : _GEN_15976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15978 = 9'hc6 == r_count_39_io_out ? io_r_198_b : _GEN_15977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15979 = 9'hc7 == r_count_39_io_out ? io_r_199_b : _GEN_15978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15980 = 9'hc8 == r_count_39_io_out ? io_r_200_b : _GEN_15979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15981 = 9'hc9 == r_count_39_io_out ? io_r_201_b : _GEN_15980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15982 = 9'hca == r_count_39_io_out ? io_r_202_b : _GEN_15981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15983 = 9'hcb == r_count_39_io_out ? io_r_203_b : _GEN_15982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15984 = 9'hcc == r_count_39_io_out ? io_r_204_b : _GEN_15983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15985 = 9'hcd == r_count_39_io_out ? io_r_205_b : _GEN_15984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15986 = 9'hce == r_count_39_io_out ? io_r_206_b : _GEN_15985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15987 = 9'hcf == r_count_39_io_out ? io_r_207_b : _GEN_15986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15988 = 9'hd0 == r_count_39_io_out ? io_r_208_b : _GEN_15987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15989 = 9'hd1 == r_count_39_io_out ? io_r_209_b : _GEN_15988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15990 = 9'hd2 == r_count_39_io_out ? io_r_210_b : _GEN_15989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15991 = 9'hd3 == r_count_39_io_out ? io_r_211_b : _GEN_15990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15992 = 9'hd4 == r_count_39_io_out ? io_r_212_b : _GEN_15991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15993 = 9'hd5 == r_count_39_io_out ? io_r_213_b : _GEN_15992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15994 = 9'hd6 == r_count_39_io_out ? io_r_214_b : _GEN_15993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15995 = 9'hd7 == r_count_39_io_out ? io_r_215_b : _GEN_15994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15996 = 9'hd8 == r_count_39_io_out ? io_r_216_b : _GEN_15995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15997 = 9'hd9 == r_count_39_io_out ? io_r_217_b : _GEN_15996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15998 = 9'hda == r_count_39_io_out ? io_r_218_b : _GEN_15997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15999 = 9'hdb == r_count_39_io_out ? io_r_219_b : _GEN_15998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16000 = 9'hdc == r_count_39_io_out ? io_r_220_b : _GEN_15999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16001 = 9'hdd == r_count_39_io_out ? io_r_221_b : _GEN_16000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16002 = 9'hde == r_count_39_io_out ? io_r_222_b : _GEN_16001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16003 = 9'hdf == r_count_39_io_out ? io_r_223_b : _GEN_16002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16004 = 9'he0 == r_count_39_io_out ? io_r_224_b : _GEN_16003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16005 = 9'he1 == r_count_39_io_out ? io_r_225_b : _GEN_16004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16006 = 9'he2 == r_count_39_io_out ? io_r_226_b : _GEN_16005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16007 = 9'he3 == r_count_39_io_out ? io_r_227_b : _GEN_16006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16008 = 9'he4 == r_count_39_io_out ? io_r_228_b : _GEN_16007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16009 = 9'he5 == r_count_39_io_out ? io_r_229_b : _GEN_16008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16010 = 9'he6 == r_count_39_io_out ? io_r_230_b : _GEN_16009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16011 = 9'he7 == r_count_39_io_out ? io_r_231_b : _GEN_16010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16012 = 9'he8 == r_count_39_io_out ? io_r_232_b : _GEN_16011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16013 = 9'he9 == r_count_39_io_out ? io_r_233_b : _GEN_16012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16014 = 9'hea == r_count_39_io_out ? io_r_234_b : _GEN_16013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16015 = 9'heb == r_count_39_io_out ? io_r_235_b : _GEN_16014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16016 = 9'hec == r_count_39_io_out ? io_r_236_b : _GEN_16015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16017 = 9'hed == r_count_39_io_out ? io_r_237_b : _GEN_16016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16018 = 9'hee == r_count_39_io_out ? io_r_238_b : _GEN_16017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16019 = 9'hef == r_count_39_io_out ? io_r_239_b : _GEN_16018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16020 = 9'hf0 == r_count_39_io_out ? io_r_240_b : _GEN_16019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16021 = 9'hf1 == r_count_39_io_out ? io_r_241_b : _GEN_16020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16022 = 9'hf2 == r_count_39_io_out ? io_r_242_b : _GEN_16021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16023 = 9'hf3 == r_count_39_io_out ? io_r_243_b : _GEN_16022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16024 = 9'hf4 == r_count_39_io_out ? io_r_244_b : _GEN_16023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16025 = 9'hf5 == r_count_39_io_out ? io_r_245_b : _GEN_16024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16026 = 9'hf6 == r_count_39_io_out ? io_r_246_b : _GEN_16025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16027 = 9'hf7 == r_count_39_io_out ? io_r_247_b : _GEN_16026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16028 = 9'hf8 == r_count_39_io_out ? io_r_248_b : _GEN_16027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16029 = 9'hf9 == r_count_39_io_out ? io_r_249_b : _GEN_16028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16030 = 9'hfa == r_count_39_io_out ? io_r_250_b : _GEN_16029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16031 = 9'hfb == r_count_39_io_out ? io_r_251_b : _GEN_16030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16032 = 9'hfc == r_count_39_io_out ? io_r_252_b : _GEN_16031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16033 = 9'hfd == r_count_39_io_out ? io_r_253_b : _GEN_16032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16034 = 9'hfe == r_count_39_io_out ? io_r_254_b : _GEN_16033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16035 = 9'hff == r_count_39_io_out ? io_r_255_b : _GEN_16034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16036 = 9'h100 == r_count_39_io_out ? io_r_256_b : _GEN_16035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16037 = 9'h101 == r_count_39_io_out ? io_r_257_b : _GEN_16036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16038 = 9'h102 == r_count_39_io_out ? io_r_258_b : _GEN_16037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16039 = 9'h103 == r_count_39_io_out ? io_r_259_b : _GEN_16038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16040 = 9'h104 == r_count_39_io_out ? io_r_260_b : _GEN_16039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16041 = 9'h105 == r_count_39_io_out ? io_r_261_b : _GEN_16040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16042 = 9'h106 == r_count_39_io_out ? io_r_262_b : _GEN_16041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16043 = 9'h107 == r_count_39_io_out ? io_r_263_b : _GEN_16042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16044 = 9'h108 == r_count_39_io_out ? io_r_264_b : _GEN_16043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16045 = 9'h109 == r_count_39_io_out ? io_r_265_b : _GEN_16044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16046 = 9'h10a == r_count_39_io_out ? io_r_266_b : _GEN_16045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16047 = 9'h10b == r_count_39_io_out ? io_r_267_b : _GEN_16046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16048 = 9'h10c == r_count_39_io_out ? io_r_268_b : _GEN_16047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16049 = 9'h10d == r_count_39_io_out ? io_r_269_b : _GEN_16048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16050 = 9'h10e == r_count_39_io_out ? io_r_270_b : _GEN_16049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16051 = 9'h10f == r_count_39_io_out ? io_r_271_b : _GEN_16050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16052 = 9'h110 == r_count_39_io_out ? io_r_272_b : _GEN_16051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16053 = 9'h111 == r_count_39_io_out ? io_r_273_b : _GEN_16052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16054 = 9'h112 == r_count_39_io_out ? io_r_274_b : _GEN_16053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16055 = 9'h113 == r_count_39_io_out ? io_r_275_b : _GEN_16054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16056 = 9'h114 == r_count_39_io_out ? io_r_276_b : _GEN_16055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16057 = 9'h115 == r_count_39_io_out ? io_r_277_b : _GEN_16056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16058 = 9'h116 == r_count_39_io_out ? io_r_278_b : _GEN_16057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16059 = 9'h117 == r_count_39_io_out ? io_r_279_b : _GEN_16058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16060 = 9'h118 == r_count_39_io_out ? io_r_280_b : _GEN_16059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16061 = 9'h119 == r_count_39_io_out ? io_r_281_b : _GEN_16060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16062 = 9'h11a == r_count_39_io_out ? io_r_282_b : _GEN_16061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16063 = 9'h11b == r_count_39_io_out ? io_r_283_b : _GEN_16062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16064 = 9'h11c == r_count_39_io_out ? io_r_284_b : _GEN_16063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16065 = 9'h11d == r_count_39_io_out ? io_r_285_b : _GEN_16064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16066 = 9'h11e == r_count_39_io_out ? io_r_286_b : _GEN_16065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16067 = 9'h11f == r_count_39_io_out ? io_r_287_b : _GEN_16066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16068 = 9'h120 == r_count_39_io_out ? io_r_288_b : _GEN_16067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16069 = 9'h121 == r_count_39_io_out ? io_r_289_b : _GEN_16068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16070 = 9'h122 == r_count_39_io_out ? io_r_290_b : _GEN_16069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16071 = 9'h123 == r_count_39_io_out ? io_r_291_b : _GEN_16070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16072 = 9'h124 == r_count_39_io_out ? io_r_292_b : _GEN_16071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16073 = 9'h125 == r_count_39_io_out ? io_r_293_b : _GEN_16072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16074 = 9'h126 == r_count_39_io_out ? io_r_294_b : _GEN_16073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16075 = 9'h127 == r_count_39_io_out ? io_r_295_b : _GEN_16074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16076 = 9'h128 == r_count_39_io_out ? io_r_296_b : _GEN_16075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16077 = 9'h129 == r_count_39_io_out ? io_r_297_b : _GEN_16076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16078 = 9'h12a == r_count_39_io_out ? io_r_298_b : _GEN_16077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16079 = 9'h12b == r_count_39_io_out ? io_r_299_b : _GEN_16078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16080 = 9'h12c == r_count_39_io_out ? io_r_300_b : _GEN_16079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16081 = 9'h12d == r_count_39_io_out ? io_r_301_b : _GEN_16080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16082 = 9'h12e == r_count_39_io_out ? io_r_302_b : _GEN_16081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16083 = 9'h12f == r_count_39_io_out ? io_r_303_b : _GEN_16082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16084 = 9'h130 == r_count_39_io_out ? io_r_304_b : _GEN_16083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16085 = 9'h131 == r_count_39_io_out ? io_r_305_b : _GEN_16084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16086 = 9'h132 == r_count_39_io_out ? io_r_306_b : _GEN_16085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16087 = 9'h133 == r_count_39_io_out ? io_r_307_b : _GEN_16086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16088 = 9'h134 == r_count_39_io_out ? io_r_308_b : _GEN_16087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16089 = 9'h135 == r_count_39_io_out ? io_r_309_b : _GEN_16088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16090 = 9'h136 == r_count_39_io_out ? io_r_310_b : _GEN_16089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16091 = 9'h137 == r_count_39_io_out ? io_r_311_b : _GEN_16090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16092 = 9'h138 == r_count_39_io_out ? io_r_312_b : _GEN_16091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16093 = 9'h139 == r_count_39_io_out ? io_r_313_b : _GEN_16092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16094 = 9'h13a == r_count_39_io_out ? io_r_314_b : _GEN_16093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16095 = 9'h13b == r_count_39_io_out ? io_r_315_b : _GEN_16094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16096 = 9'h13c == r_count_39_io_out ? io_r_316_b : _GEN_16095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16097 = 9'h13d == r_count_39_io_out ? io_r_317_b : _GEN_16096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16098 = 9'h13e == r_count_39_io_out ? io_r_318_b : _GEN_16097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16099 = 9'h13f == r_count_39_io_out ? io_r_319_b : _GEN_16098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16100 = 9'h140 == r_count_39_io_out ? io_r_320_b : _GEN_16099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16101 = 9'h141 == r_count_39_io_out ? io_r_321_b : _GEN_16100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16102 = 9'h142 == r_count_39_io_out ? io_r_322_b : _GEN_16101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16103 = 9'h143 == r_count_39_io_out ? io_r_323_b : _GEN_16102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16104 = 9'h144 == r_count_39_io_out ? io_r_324_b : _GEN_16103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16105 = 9'h145 == r_count_39_io_out ? io_r_325_b : _GEN_16104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16106 = 9'h146 == r_count_39_io_out ? io_r_326_b : _GEN_16105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16107 = 9'h147 == r_count_39_io_out ? io_r_327_b : _GEN_16106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16108 = 9'h148 == r_count_39_io_out ? io_r_328_b : _GEN_16107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16109 = 9'h149 == r_count_39_io_out ? io_r_329_b : _GEN_16108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16110 = 9'h14a == r_count_39_io_out ? io_r_330_b : _GEN_16109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16111 = 9'h14b == r_count_39_io_out ? io_r_331_b : _GEN_16110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16112 = 9'h14c == r_count_39_io_out ? io_r_332_b : _GEN_16111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16113 = 9'h14d == r_count_39_io_out ? io_r_333_b : _GEN_16112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16114 = 9'h14e == r_count_39_io_out ? io_r_334_b : _GEN_16113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16115 = 9'h14f == r_count_39_io_out ? io_r_335_b : _GEN_16114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16116 = 9'h150 == r_count_39_io_out ? io_r_336_b : _GEN_16115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16117 = 9'h151 == r_count_39_io_out ? io_r_337_b : _GEN_16116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16118 = 9'h152 == r_count_39_io_out ? io_r_338_b : _GEN_16117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16119 = 9'h153 == r_count_39_io_out ? io_r_339_b : _GEN_16118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16120 = 9'h154 == r_count_39_io_out ? io_r_340_b : _GEN_16119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16121 = 9'h155 == r_count_39_io_out ? io_r_341_b : _GEN_16120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16122 = 9'h156 == r_count_39_io_out ? io_r_342_b : _GEN_16121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16123 = 9'h157 == r_count_39_io_out ? io_r_343_b : _GEN_16122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16124 = 9'h158 == r_count_39_io_out ? io_r_344_b : _GEN_16123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16125 = 9'h159 == r_count_39_io_out ? io_r_345_b : _GEN_16124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16126 = 9'h15a == r_count_39_io_out ? io_r_346_b : _GEN_16125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16127 = 9'h15b == r_count_39_io_out ? io_r_347_b : _GEN_16126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16128 = 9'h15c == r_count_39_io_out ? io_r_348_b : _GEN_16127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16129 = 9'h15d == r_count_39_io_out ? io_r_349_b : _GEN_16128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16130 = 9'h15e == r_count_39_io_out ? io_r_350_b : _GEN_16129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16131 = 9'h15f == r_count_39_io_out ? io_r_351_b : _GEN_16130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16132 = 9'h160 == r_count_39_io_out ? io_r_352_b : _GEN_16131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16133 = 9'h161 == r_count_39_io_out ? io_r_353_b : _GEN_16132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16134 = 9'h162 == r_count_39_io_out ? io_r_354_b : _GEN_16133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16135 = 9'h163 == r_count_39_io_out ? io_r_355_b : _GEN_16134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16136 = 9'h164 == r_count_39_io_out ? io_r_356_b : _GEN_16135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16137 = 9'h165 == r_count_39_io_out ? io_r_357_b : _GEN_16136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16138 = 9'h166 == r_count_39_io_out ? io_r_358_b : _GEN_16137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16139 = 9'h167 == r_count_39_io_out ? io_r_359_b : _GEN_16138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16140 = 9'h168 == r_count_39_io_out ? io_r_360_b : _GEN_16139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16141 = 9'h169 == r_count_39_io_out ? io_r_361_b : _GEN_16140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16142 = 9'h16a == r_count_39_io_out ? io_r_362_b : _GEN_16141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16143 = 9'h16b == r_count_39_io_out ? io_r_363_b : _GEN_16142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16144 = 9'h16c == r_count_39_io_out ? io_r_364_b : _GEN_16143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16145 = 9'h16d == r_count_39_io_out ? io_r_365_b : _GEN_16144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16146 = 9'h16e == r_count_39_io_out ? io_r_366_b : _GEN_16145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16147 = 9'h16f == r_count_39_io_out ? io_r_367_b : _GEN_16146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16148 = 9'h170 == r_count_39_io_out ? io_r_368_b : _GEN_16147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16149 = 9'h171 == r_count_39_io_out ? io_r_369_b : _GEN_16148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16150 = 9'h172 == r_count_39_io_out ? io_r_370_b : _GEN_16149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16151 = 9'h173 == r_count_39_io_out ? io_r_371_b : _GEN_16150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16152 = 9'h174 == r_count_39_io_out ? io_r_372_b : _GEN_16151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16153 = 9'h175 == r_count_39_io_out ? io_r_373_b : _GEN_16152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16154 = 9'h176 == r_count_39_io_out ? io_r_374_b : _GEN_16153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16155 = 9'h177 == r_count_39_io_out ? io_r_375_b : _GEN_16154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16156 = 9'h178 == r_count_39_io_out ? io_r_376_b : _GEN_16155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16157 = 9'h179 == r_count_39_io_out ? io_r_377_b : _GEN_16156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16158 = 9'h17a == r_count_39_io_out ? io_r_378_b : _GEN_16157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16159 = 9'h17b == r_count_39_io_out ? io_r_379_b : _GEN_16158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16160 = 9'h17c == r_count_39_io_out ? io_r_380_b : _GEN_16159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16161 = 9'h17d == r_count_39_io_out ? io_r_381_b : _GEN_16160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16162 = 9'h17e == r_count_39_io_out ? io_r_382_b : _GEN_16161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16163 = 9'h17f == r_count_39_io_out ? io_r_383_b : _GEN_16162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16164 = 9'h180 == r_count_39_io_out ? io_r_384_b : _GEN_16163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16165 = 9'h181 == r_count_39_io_out ? io_r_385_b : _GEN_16164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16166 = 9'h182 == r_count_39_io_out ? io_r_386_b : _GEN_16165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16167 = 9'h183 == r_count_39_io_out ? io_r_387_b : _GEN_16166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16168 = 9'h184 == r_count_39_io_out ? io_r_388_b : _GEN_16167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16169 = 9'h185 == r_count_39_io_out ? io_r_389_b : _GEN_16168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16170 = 9'h186 == r_count_39_io_out ? io_r_390_b : _GEN_16169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16171 = 9'h187 == r_count_39_io_out ? io_r_391_b : _GEN_16170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16172 = 9'h188 == r_count_39_io_out ? io_r_392_b : _GEN_16171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16173 = 9'h189 == r_count_39_io_out ? io_r_393_b : _GEN_16172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16174 = 9'h18a == r_count_39_io_out ? io_r_394_b : _GEN_16173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16175 = 9'h18b == r_count_39_io_out ? io_r_395_b : _GEN_16174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16176 = 9'h18c == r_count_39_io_out ? io_r_396_b : _GEN_16175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16177 = 9'h18d == r_count_39_io_out ? io_r_397_b : _GEN_16176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16178 = 9'h18e == r_count_39_io_out ? io_r_398_b : _GEN_16177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16181 = 9'h1 == r_count_40_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16182 = 9'h2 == r_count_40_io_out ? io_r_2_b : _GEN_16181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16183 = 9'h3 == r_count_40_io_out ? io_r_3_b : _GEN_16182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16184 = 9'h4 == r_count_40_io_out ? io_r_4_b : _GEN_16183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16185 = 9'h5 == r_count_40_io_out ? io_r_5_b : _GEN_16184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16186 = 9'h6 == r_count_40_io_out ? io_r_6_b : _GEN_16185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16187 = 9'h7 == r_count_40_io_out ? io_r_7_b : _GEN_16186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16188 = 9'h8 == r_count_40_io_out ? io_r_8_b : _GEN_16187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16189 = 9'h9 == r_count_40_io_out ? io_r_9_b : _GEN_16188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16190 = 9'ha == r_count_40_io_out ? io_r_10_b : _GEN_16189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16191 = 9'hb == r_count_40_io_out ? io_r_11_b : _GEN_16190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16192 = 9'hc == r_count_40_io_out ? io_r_12_b : _GEN_16191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16193 = 9'hd == r_count_40_io_out ? io_r_13_b : _GEN_16192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16194 = 9'he == r_count_40_io_out ? io_r_14_b : _GEN_16193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16195 = 9'hf == r_count_40_io_out ? io_r_15_b : _GEN_16194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16196 = 9'h10 == r_count_40_io_out ? io_r_16_b : _GEN_16195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16197 = 9'h11 == r_count_40_io_out ? io_r_17_b : _GEN_16196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16198 = 9'h12 == r_count_40_io_out ? io_r_18_b : _GEN_16197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16199 = 9'h13 == r_count_40_io_out ? io_r_19_b : _GEN_16198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16200 = 9'h14 == r_count_40_io_out ? io_r_20_b : _GEN_16199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16201 = 9'h15 == r_count_40_io_out ? io_r_21_b : _GEN_16200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16202 = 9'h16 == r_count_40_io_out ? io_r_22_b : _GEN_16201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16203 = 9'h17 == r_count_40_io_out ? io_r_23_b : _GEN_16202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16204 = 9'h18 == r_count_40_io_out ? io_r_24_b : _GEN_16203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16205 = 9'h19 == r_count_40_io_out ? io_r_25_b : _GEN_16204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16206 = 9'h1a == r_count_40_io_out ? io_r_26_b : _GEN_16205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16207 = 9'h1b == r_count_40_io_out ? io_r_27_b : _GEN_16206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16208 = 9'h1c == r_count_40_io_out ? io_r_28_b : _GEN_16207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16209 = 9'h1d == r_count_40_io_out ? io_r_29_b : _GEN_16208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16210 = 9'h1e == r_count_40_io_out ? io_r_30_b : _GEN_16209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16211 = 9'h1f == r_count_40_io_out ? io_r_31_b : _GEN_16210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16212 = 9'h20 == r_count_40_io_out ? io_r_32_b : _GEN_16211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16213 = 9'h21 == r_count_40_io_out ? io_r_33_b : _GEN_16212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16214 = 9'h22 == r_count_40_io_out ? io_r_34_b : _GEN_16213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16215 = 9'h23 == r_count_40_io_out ? io_r_35_b : _GEN_16214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16216 = 9'h24 == r_count_40_io_out ? io_r_36_b : _GEN_16215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16217 = 9'h25 == r_count_40_io_out ? io_r_37_b : _GEN_16216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16218 = 9'h26 == r_count_40_io_out ? io_r_38_b : _GEN_16217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16219 = 9'h27 == r_count_40_io_out ? io_r_39_b : _GEN_16218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16220 = 9'h28 == r_count_40_io_out ? io_r_40_b : _GEN_16219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16221 = 9'h29 == r_count_40_io_out ? io_r_41_b : _GEN_16220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16222 = 9'h2a == r_count_40_io_out ? io_r_42_b : _GEN_16221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16223 = 9'h2b == r_count_40_io_out ? io_r_43_b : _GEN_16222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16224 = 9'h2c == r_count_40_io_out ? io_r_44_b : _GEN_16223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16225 = 9'h2d == r_count_40_io_out ? io_r_45_b : _GEN_16224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16226 = 9'h2e == r_count_40_io_out ? io_r_46_b : _GEN_16225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16227 = 9'h2f == r_count_40_io_out ? io_r_47_b : _GEN_16226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16228 = 9'h30 == r_count_40_io_out ? io_r_48_b : _GEN_16227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16229 = 9'h31 == r_count_40_io_out ? io_r_49_b : _GEN_16228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16230 = 9'h32 == r_count_40_io_out ? io_r_50_b : _GEN_16229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16231 = 9'h33 == r_count_40_io_out ? io_r_51_b : _GEN_16230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16232 = 9'h34 == r_count_40_io_out ? io_r_52_b : _GEN_16231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16233 = 9'h35 == r_count_40_io_out ? io_r_53_b : _GEN_16232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16234 = 9'h36 == r_count_40_io_out ? io_r_54_b : _GEN_16233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16235 = 9'h37 == r_count_40_io_out ? io_r_55_b : _GEN_16234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16236 = 9'h38 == r_count_40_io_out ? io_r_56_b : _GEN_16235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16237 = 9'h39 == r_count_40_io_out ? io_r_57_b : _GEN_16236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16238 = 9'h3a == r_count_40_io_out ? io_r_58_b : _GEN_16237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16239 = 9'h3b == r_count_40_io_out ? io_r_59_b : _GEN_16238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16240 = 9'h3c == r_count_40_io_out ? io_r_60_b : _GEN_16239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16241 = 9'h3d == r_count_40_io_out ? io_r_61_b : _GEN_16240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16242 = 9'h3e == r_count_40_io_out ? io_r_62_b : _GEN_16241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16243 = 9'h3f == r_count_40_io_out ? io_r_63_b : _GEN_16242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16244 = 9'h40 == r_count_40_io_out ? io_r_64_b : _GEN_16243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16245 = 9'h41 == r_count_40_io_out ? io_r_65_b : _GEN_16244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16246 = 9'h42 == r_count_40_io_out ? io_r_66_b : _GEN_16245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16247 = 9'h43 == r_count_40_io_out ? io_r_67_b : _GEN_16246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16248 = 9'h44 == r_count_40_io_out ? io_r_68_b : _GEN_16247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16249 = 9'h45 == r_count_40_io_out ? io_r_69_b : _GEN_16248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16250 = 9'h46 == r_count_40_io_out ? io_r_70_b : _GEN_16249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16251 = 9'h47 == r_count_40_io_out ? io_r_71_b : _GEN_16250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16252 = 9'h48 == r_count_40_io_out ? io_r_72_b : _GEN_16251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16253 = 9'h49 == r_count_40_io_out ? io_r_73_b : _GEN_16252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16254 = 9'h4a == r_count_40_io_out ? io_r_74_b : _GEN_16253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16255 = 9'h4b == r_count_40_io_out ? io_r_75_b : _GEN_16254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16256 = 9'h4c == r_count_40_io_out ? io_r_76_b : _GEN_16255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16257 = 9'h4d == r_count_40_io_out ? io_r_77_b : _GEN_16256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16258 = 9'h4e == r_count_40_io_out ? io_r_78_b : _GEN_16257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16259 = 9'h4f == r_count_40_io_out ? io_r_79_b : _GEN_16258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16260 = 9'h50 == r_count_40_io_out ? io_r_80_b : _GEN_16259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16261 = 9'h51 == r_count_40_io_out ? io_r_81_b : _GEN_16260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16262 = 9'h52 == r_count_40_io_out ? io_r_82_b : _GEN_16261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16263 = 9'h53 == r_count_40_io_out ? io_r_83_b : _GEN_16262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16264 = 9'h54 == r_count_40_io_out ? io_r_84_b : _GEN_16263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16265 = 9'h55 == r_count_40_io_out ? io_r_85_b : _GEN_16264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16266 = 9'h56 == r_count_40_io_out ? io_r_86_b : _GEN_16265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16267 = 9'h57 == r_count_40_io_out ? io_r_87_b : _GEN_16266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16268 = 9'h58 == r_count_40_io_out ? io_r_88_b : _GEN_16267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16269 = 9'h59 == r_count_40_io_out ? io_r_89_b : _GEN_16268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16270 = 9'h5a == r_count_40_io_out ? io_r_90_b : _GEN_16269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16271 = 9'h5b == r_count_40_io_out ? io_r_91_b : _GEN_16270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16272 = 9'h5c == r_count_40_io_out ? io_r_92_b : _GEN_16271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16273 = 9'h5d == r_count_40_io_out ? io_r_93_b : _GEN_16272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16274 = 9'h5e == r_count_40_io_out ? io_r_94_b : _GEN_16273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16275 = 9'h5f == r_count_40_io_out ? io_r_95_b : _GEN_16274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16276 = 9'h60 == r_count_40_io_out ? io_r_96_b : _GEN_16275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16277 = 9'h61 == r_count_40_io_out ? io_r_97_b : _GEN_16276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16278 = 9'h62 == r_count_40_io_out ? io_r_98_b : _GEN_16277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16279 = 9'h63 == r_count_40_io_out ? io_r_99_b : _GEN_16278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16280 = 9'h64 == r_count_40_io_out ? io_r_100_b : _GEN_16279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16281 = 9'h65 == r_count_40_io_out ? io_r_101_b : _GEN_16280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16282 = 9'h66 == r_count_40_io_out ? io_r_102_b : _GEN_16281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16283 = 9'h67 == r_count_40_io_out ? io_r_103_b : _GEN_16282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16284 = 9'h68 == r_count_40_io_out ? io_r_104_b : _GEN_16283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16285 = 9'h69 == r_count_40_io_out ? io_r_105_b : _GEN_16284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16286 = 9'h6a == r_count_40_io_out ? io_r_106_b : _GEN_16285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16287 = 9'h6b == r_count_40_io_out ? io_r_107_b : _GEN_16286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16288 = 9'h6c == r_count_40_io_out ? io_r_108_b : _GEN_16287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16289 = 9'h6d == r_count_40_io_out ? io_r_109_b : _GEN_16288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16290 = 9'h6e == r_count_40_io_out ? io_r_110_b : _GEN_16289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16291 = 9'h6f == r_count_40_io_out ? io_r_111_b : _GEN_16290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16292 = 9'h70 == r_count_40_io_out ? io_r_112_b : _GEN_16291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16293 = 9'h71 == r_count_40_io_out ? io_r_113_b : _GEN_16292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16294 = 9'h72 == r_count_40_io_out ? io_r_114_b : _GEN_16293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16295 = 9'h73 == r_count_40_io_out ? io_r_115_b : _GEN_16294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16296 = 9'h74 == r_count_40_io_out ? io_r_116_b : _GEN_16295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16297 = 9'h75 == r_count_40_io_out ? io_r_117_b : _GEN_16296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16298 = 9'h76 == r_count_40_io_out ? io_r_118_b : _GEN_16297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16299 = 9'h77 == r_count_40_io_out ? io_r_119_b : _GEN_16298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16300 = 9'h78 == r_count_40_io_out ? io_r_120_b : _GEN_16299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16301 = 9'h79 == r_count_40_io_out ? io_r_121_b : _GEN_16300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16302 = 9'h7a == r_count_40_io_out ? io_r_122_b : _GEN_16301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16303 = 9'h7b == r_count_40_io_out ? io_r_123_b : _GEN_16302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16304 = 9'h7c == r_count_40_io_out ? io_r_124_b : _GEN_16303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16305 = 9'h7d == r_count_40_io_out ? io_r_125_b : _GEN_16304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16306 = 9'h7e == r_count_40_io_out ? io_r_126_b : _GEN_16305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16307 = 9'h7f == r_count_40_io_out ? io_r_127_b : _GEN_16306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16308 = 9'h80 == r_count_40_io_out ? io_r_128_b : _GEN_16307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16309 = 9'h81 == r_count_40_io_out ? io_r_129_b : _GEN_16308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16310 = 9'h82 == r_count_40_io_out ? io_r_130_b : _GEN_16309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16311 = 9'h83 == r_count_40_io_out ? io_r_131_b : _GEN_16310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16312 = 9'h84 == r_count_40_io_out ? io_r_132_b : _GEN_16311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16313 = 9'h85 == r_count_40_io_out ? io_r_133_b : _GEN_16312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16314 = 9'h86 == r_count_40_io_out ? io_r_134_b : _GEN_16313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16315 = 9'h87 == r_count_40_io_out ? io_r_135_b : _GEN_16314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16316 = 9'h88 == r_count_40_io_out ? io_r_136_b : _GEN_16315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16317 = 9'h89 == r_count_40_io_out ? io_r_137_b : _GEN_16316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16318 = 9'h8a == r_count_40_io_out ? io_r_138_b : _GEN_16317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16319 = 9'h8b == r_count_40_io_out ? io_r_139_b : _GEN_16318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16320 = 9'h8c == r_count_40_io_out ? io_r_140_b : _GEN_16319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16321 = 9'h8d == r_count_40_io_out ? io_r_141_b : _GEN_16320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16322 = 9'h8e == r_count_40_io_out ? io_r_142_b : _GEN_16321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16323 = 9'h8f == r_count_40_io_out ? io_r_143_b : _GEN_16322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16324 = 9'h90 == r_count_40_io_out ? io_r_144_b : _GEN_16323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16325 = 9'h91 == r_count_40_io_out ? io_r_145_b : _GEN_16324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16326 = 9'h92 == r_count_40_io_out ? io_r_146_b : _GEN_16325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16327 = 9'h93 == r_count_40_io_out ? io_r_147_b : _GEN_16326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16328 = 9'h94 == r_count_40_io_out ? io_r_148_b : _GEN_16327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16329 = 9'h95 == r_count_40_io_out ? io_r_149_b : _GEN_16328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16330 = 9'h96 == r_count_40_io_out ? io_r_150_b : _GEN_16329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16331 = 9'h97 == r_count_40_io_out ? io_r_151_b : _GEN_16330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16332 = 9'h98 == r_count_40_io_out ? io_r_152_b : _GEN_16331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16333 = 9'h99 == r_count_40_io_out ? io_r_153_b : _GEN_16332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16334 = 9'h9a == r_count_40_io_out ? io_r_154_b : _GEN_16333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16335 = 9'h9b == r_count_40_io_out ? io_r_155_b : _GEN_16334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16336 = 9'h9c == r_count_40_io_out ? io_r_156_b : _GEN_16335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16337 = 9'h9d == r_count_40_io_out ? io_r_157_b : _GEN_16336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16338 = 9'h9e == r_count_40_io_out ? io_r_158_b : _GEN_16337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16339 = 9'h9f == r_count_40_io_out ? io_r_159_b : _GEN_16338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16340 = 9'ha0 == r_count_40_io_out ? io_r_160_b : _GEN_16339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16341 = 9'ha1 == r_count_40_io_out ? io_r_161_b : _GEN_16340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16342 = 9'ha2 == r_count_40_io_out ? io_r_162_b : _GEN_16341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16343 = 9'ha3 == r_count_40_io_out ? io_r_163_b : _GEN_16342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16344 = 9'ha4 == r_count_40_io_out ? io_r_164_b : _GEN_16343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16345 = 9'ha5 == r_count_40_io_out ? io_r_165_b : _GEN_16344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16346 = 9'ha6 == r_count_40_io_out ? io_r_166_b : _GEN_16345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16347 = 9'ha7 == r_count_40_io_out ? io_r_167_b : _GEN_16346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16348 = 9'ha8 == r_count_40_io_out ? io_r_168_b : _GEN_16347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16349 = 9'ha9 == r_count_40_io_out ? io_r_169_b : _GEN_16348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16350 = 9'haa == r_count_40_io_out ? io_r_170_b : _GEN_16349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16351 = 9'hab == r_count_40_io_out ? io_r_171_b : _GEN_16350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16352 = 9'hac == r_count_40_io_out ? io_r_172_b : _GEN_16351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16353 = 9'had == r_count_40_io_out ? io_r_173_b : _GEN_16352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16354 = 9'hae == r_count_40_io_out ? io_r_174_b : _GEN_16353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16355 = 9'haf == r_count_40_io_out ? io_r_175_b : _GEN_16354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16356 = 9'hb0 == r_count_40_io_out ? io_r_176_b : _GEN_16355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16357 = 9'hb1 == r_count_40_io_out ? io_r_177_b : _GEN_16356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16358 = 9'hb2 == r_count_40_io_out ? io_r_178_b : _GEN_16357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16359 = 9'hb3 == r_count_40_io_out ? io_r_179_b : _GEN_16358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16360 = 9'hb4 == r_count_40_io_out ? io_r_180_b : _GEN_16359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16361 = 9'hb5 == r_count_40_io_out ? io_r_181_b : _GEN_16360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16362 = 9'hb6 == r_count_40_io_out ? io_r_182_b : _GEN_16361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16363 = 9'hb7 == r_count_40_io_out ? io_r_183_b : _GEN_16362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16364 = 9'hb8 == r_count_40_io_out ? io_r_184_b : _GEN_16363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16365 = 9'hb9 == r_count_40_io_out ? io_r_185_b : _GEN_16364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16366 = 9'hba == r_count_40_io_out ? io_r_186_b : _GEN_16365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16367 = 9'hbb == r_count_40_io_out ? io_r_187_b : _GEN_16366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16368 = 9'hbc == r_count_40_io_out ? io_r_188_b : _GEN_16367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16369 = 9'hbd == r_count_40_io_out ? io_r_189_b : _GEN_16368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16370 = 9'hbe == r_count_40_io_out ? io_r_190_b : _GEN_16369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16371 = 9'hbf == r_count_40_io_out ? io_r_191_b : _GEN_16370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16372 = 9'hc0 == r_count_40_io_out ? io_r_192_b : _GEN_16371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16373 = 9'hc1 == r_count_40_io_out ? io_r_193_b : _GEN_16372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16374 = 9'hc2 == r_count_40_io_out ? io_r_194_b : _GEN_16373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16375 = 9'hc3 == r_count_40_io_out ? io_r_195_b : _GEN_16374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16376 = 9'hc4 == r_count_40_io_out ? io_r_196_b : _GEN_16375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16377 = 9'hc5 == r_count_40_io_out ? io_r_197_b : _GEN_16376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16378 = 9'hc6 == r_count_40_io_out ? io_r_198_b : _GEN_16377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16379 = 9'hc7 == r_count_40_io_out ? io_r_199_b : _GEN_16378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16380 = 9'hc8 == r_count_40_io_out ? io_r_200_b : _GEN_16379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16381 = 9'hc9 == r_count_40_io_out ? io_r_201_b : _GEN_16380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16382 = 9'hca == r_count_40_io_out ? io_r_202_b : _GEN_16381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16383 = 9'hcb == r_count_40_io_out ? io_r_203_b : _GEN_16382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16384 = 9'hcc == r_count_40_io_out ? io_r_204_b : _GEN_16383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16385 = 9'hcd == r_count_40_io_out ? io_r_205_b : _GEN_16384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16386 = 9'hce == r_count_40_io_out ? io_r_206_b : _GEN_16385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16387 = 9'hcf == r_count_40_io_out ? io_r_207_b : _GEN_16386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16388 = 9'hd0 == r_count_40_io_out ? io_r_208_b : _GEN_16387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16389 = 9'hd1 == r_count_40_io_out ? io_r_209_b : _GEN_16388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16390 = 9'hd2 == r_count_40_io_out ? io_r_210_b : _GEN_16389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16391 = 9'hd3 == r_count_40_io_out ? io_r_211_b : _GEN_16390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16392 = 9'hd4 == r_count_40_io_out ? io_r_212_b : _GEN_16391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16393 = 9'hd5 == r_count_40_io_out ? io_r_213_b : _GEN_16392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16394 = 9'hd6 == r_count_40_io_out ? io_r_214_b : _GEN_16393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16395 = 9'hd7 == r_count_40_io_out ? io_r_215_b : _GEN_16394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16396 = 9'hd8 == r_count_40_io_out ? io_r_216_b : _GEN_16395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16397 = 9'hd9 == r_count_40_io_out ? io_r_217_b : _GEN_16396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16398 = 9'hda == r_count_40_io_out ? io_r_218_b : _GEN_16397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16399 = 9'hdb == r_count_40_io_out ? io_r_219_b : _GEN_16398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16400 = 9'hdc == r_count_40_io_out ? io_r_220_b : _GEN_16399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16401 = 9'hdd == r_count_40_io_out ? io_r_221_b : _GEN_16400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16402 = 9'hde == r_count_40_io_out ? io_r_222_b : _GEN_16401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16403 = 9'hdf == r_count_40_io_out ? io_r_223_b : _GEN_16402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16404 = 9'he0 == r_count_40_io_out ? io_r_224_b : _GEN_16403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16405 = 9'he1 == r_count_40_io_out ? io_r_225_b : _GEN_16404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16406 = 9'he2 == r_count_40_io_out ? io_r_226_b : _GEN_16405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16407 = 9'he3 == r_count_40_io_out ? io_r_227_b : _GEN_16406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16408 = 9'he4 == r_count_40_io_out ? io_r_228_b : _GEN_16407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16409 = 9'he5 == r_count_40_io_out ? io_r_229_b : _GEN_16408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16410 = 9'he6 == r_count_40_io_out ? io_r_230_b : _GEN_16409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16411 = 9'he7 == r_count_40_io_out ? io_r_231_b : _GEN_16410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16412 = 9'he8 == r_count_40_io_out ? io_r_232_b : _GEN_16411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16413 = 9'he9 == r_count_40_io_out ? io_r_233_b : _GEN_16412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16414 = 9'hea == r_count_40_io_out ? io_r_234_b : _GEN_16413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16415 = 9'heb == r_count_40_io_out ? io_r_235_b : _GEN_16414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16416 = 9'hec == r_count_40_io_out ? io_r_236_b : _GEN_16415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16417 = 9'hed == r_count_40_io_out ? io_r_237_b : _GEN_16416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16418 = 9'hee == r_count_40_io_out ? io_r_238_b : _GEN_16417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16419 = 9'hef == r_count_40_io_out ? io_r_239_b : _GEN_16418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16420 = 9'hf0 == r_count_40_io_out ? io_r_240_b : _GEN_16419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16421 = 9'hf1 == r_count_40_io_out ? io_r_241_b : _GEN_16420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16422 = 9'hf2 == r_count_40_io_out ? io_r_242_b : _GEN_16421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16423 = 9'hf3 == r_count_40_io_out ? io_r_243_b : _GEN_16422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16424 = 9'hf4 == r_count_40_io_out ? io_r_244_b : _GEN_16423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16425 = 9'hf5 == r_count_40_io_out ? io_r_245_b : _GEN_16424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16426 = 9'hf6 == r_count_40_io_out ? io_r_246_b : _GEN_16425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16427 = 9'hf7 == r_count_40_io_out ? io_r_247_b : _GEN_16426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16428 = 9'hf8 == r_count_40_io_out ? io_r_248_b : _GEN_16427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16429 = 9'hf9 == r_count_40_io_out ? io_r_249_b : _GEN_16428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16430 = 9'hfa == r_count_40_io_out ? io_r_250_b : _GEN_16429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16431 = 9'hfb == r_count_40_io_out ? io_r_251_b : _GEN_16430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16432 = 9'hfc == r_count_40_io_out ? io_r_252_b : _GEN_16431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16433 = 9'hfd == r_count_40_io_out ? io_r_253_b : _GEN_16432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16434 = 9'hfe == r_count_40_io_out ? io_r_254_b : _GEN_16433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16435 = 9'hff == r_count_40_io_out ? io_r_255_b : _GEN_16434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16436 = 9'h100 == r_count_40_io_out ? io_r_256_b : _GEN_16435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16437 = 9'h101 == r_count_40_io_out ? io_r_257_b : _GEN_16436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16438 = 9'h102 == r_count_40_io_out ? io_r_258_b : _GEN_16437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16439 = 9'h103 == r_count_40_io_out ? io_r_259_b : _GEN_16438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16440 = 9'h104 == r_count_40_io_out ? io_r_260_b : _GEN_16439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16441 = 9'h105 == r_count_40_io_out ? io_r_261_b : _GEN_16440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16442 = 9'h106 == r_count_40_io_out ? io_r_262_b : _GEN_16441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16443 = 9'h107 == r_count_40_io_out ? io_r_263_b : _GEN_16442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16444 = 9'h108 == r_count_40_io_out ? io_r_264_b : _GEN_16443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16445 = 9'h109 == r_count_40_io_out ? io_r_265_b : _GEN_16444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16446 = 9'h10a == r_count_40_io_out ? io_r_266_b : _GEN_16445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16447 = 9'h10b == r_count_40_io_out ? io_r_267_b : _GEN_16446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16448 = 9'h10c == r_count_40_io_out ? io_r_268_b : _GEN_16447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16449 = 9'h10d == r_count_40_io_out ? io_r_269_b : _GEN_16448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16450 = 9'h10e == r_count_40_io_out ? io_r_270_b : _GEN_16449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16451 = 9'h10f == r_count_40_io_out ? io_r_271_b : _GEN_16450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16452 = 9'h110 == r_count_40_io_out ? io_r_272_b : _GEN_16451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16453 = 9'h111 == r_count_40_io_out ? io_r_273_b : _GEN_16452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16454 = 9'h112 == r_count_40_io_out ? io_r_274_b : _GEN_16453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16455 = 9'h113 == r_count_40_io_out ? io_r_275_b : _GEN_16454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16456 = 9'h114 == r_count_40_io_out ? io_r_276_b : _GEN_16455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16457 = 9'h115 == r_count_40_io_out ? io_r_277_b : _GEN_16456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16458 = 9'h116 == r_count_40_io_out ? io_r_278_b : _GEN_16457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16459 = 9'h117 == r_count_40_io_out ? io_r_279_b : _GEN_16458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16460 = 9'h118 == r_count_40_io_out ? io_r_280_b : _GEN_16459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16461 = 9'h119 == r_count_40_io_out ? io_r_281_b : _GEN_16460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16462 = 9'h11a == r_count_40_io_out ? io_r_282_b : _GEN_16461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16463 = 9'h11b == r_count_40_io_out ? io_r_283_b : _GEN_16462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16464 = 9'h11c == r_count_40_io_out ? io_r_284_b : _GEN_16463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16465 = 9'h11d == r_count_40_io_out ? io_r_285_b : _GEN_16464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16466 = 9'h11e == r_count_40_io_out ? io_r_286_b : _GEN_16465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16467 = 9'h11f == r_count_40_io_out ? io_r_287_b : _GEN_16466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16468 = 9'h120 == r_count_40_io_out ? io_r_288_b : _GEN_16467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16469 = 9'h121 == r_count_40_io_out ? io_r_289_b : _GEN_16468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16470 = 9'h122 == r_count_40_io_out ? io_r_290_b : _GEN_16469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16471 = 9'h123 == r_count_40_io_out ? io_r_291_b : _GEN_16470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16472 = 9'h124 == r_count_40_io_out ? io_r_292_b : _GEN_16471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16473 = 9'h125 == r_count_40_io_out ? io_r_293_b : _GEN_16472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16474 = 9'h126 == r_count_40_io_out ? io_r_294_b : _GEN_16473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16475 = 9'h127 == r_count_40_io_out ? io_r_295_b : _GEN_16474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16476 = 9'h128 == r_count_40_io_out ? io_r_296_b : _GEN_16475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16477 = 9'h129 == r_count_40_io_out ? io_r_297_b : _GEN_16476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16478 = 9'h12a == r_count_40_io_out ? io_r_298_b : _GEN_16477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16479 = 9'h12b == r_count_40_io_out ? io_r_299_b : _GEN_16478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16480 = 9'h12c == r_count_40_io_out ? io_r_300_b : _GEN_16479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16481 = 9'h12d == r_count_40_io_out ? io_r_301_b : _GEN_16480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16482 = 9'h12e == r_count_40_io_out ? io_r_302_b : _GEN_16481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16483 = 9'h12f == r_count_40_io_out ? io_r_303_b : _GEN_16482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16484 = 9'h130 == r_count_40_io_out ? io_r_304_b : _GEN_16483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16485 = 9'h131 == r_count_40_io_out ? io_r_305_b : _GEN_16484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16486 = 9'h132 == r_count_40_io_out ? io_r_306_b : _GEN_16485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16487 = 9'h133 == r_count_40_io_out ? io_r_307_b : _GEN_16486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16488 = 9'h134 == r_count_40_io_out ? io_r_308_b : _GEN_16487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16489 = 9'h135 == r_count_40_io_out ? io_r_309_b : _GEN_16488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16490 = 9'h136 == r_count_40_io_out ? io_r_310_b : _GEN_16489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16491 = 9'h137 == r_count_40_io_out ? io_r_311_b : _GEN_16490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16492 = 9'h138 == r_count_40_io_out ? io_r_312_b : _GEN_16491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16493 = 9'h139 == r_count_40_io_out ? io_r_313_b : _GEN_16492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16494 = 9'h13a == r_count_40_io_out ? io_r_314_b : _GEN_16493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16495 = 9'h13b == r_count_40_io_out ? io_r_315_b : _GEN_16494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16496 = 9'h13c == r_count_40_io_out ? io_r_316_b : _GEN_16495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16497 = 9'h13d == r_count_40_io_out ? io_r_317_b : _GEN_16496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16498 = 9'h13e == r_count_40_io_out ? io_r_318_b : _GEN_16497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16499 = 9'h13f == r_count_40_io_out ? io_r_319_b : _GEN_16498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16500 = 9'h140 == r_count_40_io_out ? io_r_320_b : _GEN_16499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16501 = 9'h141 == r_count_40_io_out ? io_r_321_b : _GEN_16500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16502 = 9'h142 == r_count_40_io_out ? io_r_322_b : _GEN_16501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16503 = 9'h143 == r_count_40_io_out ? io_r_323_b : _GEN_16502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16504 = 9'h144 == r_count_40_io_out ? io_r_324_b : _GEN_16503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16505 = 9'h145 == r_count_40_io_out ? io_r_325_b : _GEN_16504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16506 = 9'h146 == r_count_40_io_out ? io_r_326_b : _GEN_16505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16507 = 9'h147 == r_count_40_io_out ? io_r_327_b : _GEN_16506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16508 = 9'h148 == r_count_40_io_out ? io_r_328_b : _GEN_16507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16509 = 9'h149 == r_count_40_io_out ? io_r_329_b : _GEN_16508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16510 = 9'h14a == r_count_40_io_out ? io_r_330_b : _GEN_16509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16511 = 9'h14b == r_count_40_io_out ? io_r_331_b : _GEN_16510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16512 = 9'h14c == r_count_40_io_out ? io_r_332_b : _GEN_16511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16513 = 9'h14d == r_count_40_io_out ? io_r_333_b : _GEN_16512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16514 = 9'h14e == r_count_40_io_out ? io_r_334_b : _GEN_16513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16515 = 9'h14f == r_count_40_io_out ? io_r_335_b : _GEN_16514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16516 = 9'h150 == r_count_40_io_out ? io_r_336_b : _GEN_16515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16517 = 9'h151 == r_count_40_io_out ? io_r_337_b : _GEN_16516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16518 = 9'h152 == r_count_40_io_out ? io_r_338_b : _GEN_16517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16519 = 9'h153 == r_count_40_io_out ? io_r_339_b : _GEN_16518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16520 = 9'h154 == r_count_40_io_out ? io_r_340_b : _GEN_16519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16521 = 9'h155 == r_count_40_io_out ? io_r_341_b : _GEN_16520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16522 = 9'h156 == r_count_40_io_out ? io_r_342_b : _GEN_16521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16523 = 9'h157 == r_count_40_io_out ? io_r_343_b : _GEN_16522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16524 = 9'h158 == r_count_40_io_out ? io_r_344_b : _GEN_16523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16525 = 9'h159 == r_count_40_io_out ? io_r_345_b : _GEN_16524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16526 = 9'h15a == r_count_40_io_out ? io_r_346_b : _GEN_16525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16527 = 9'h15b == r_count_40_io_out ? io_r_347_b : _GEN_16526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16528 = 9'h15c == r_count_40_io_out ? io_r_348_b : _GEN_16527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16529 = 9'h15d == r_count_40_io_out ? io_r_349_b : _GEN_16528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16530 = 9'h15e == r_count_40_io_out ? io_r_350_b : _GEN_16529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16531 = 9'h15f == r_count_40_io_out ? io_r_351_b : _GEN_16530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16532 = 9'h160 == r_count_40_io_out ? io_r_352_b : _GEN_16531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16533 = 9'h161 == r_count_40_io_out ? io_r_353_b : _GEN_16532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16534 = 9'h162 == r_count_40_io_out ? io_r_354_b : _GEN_16533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16535 = 9'h163 == r_count_40_io_out ? io_r_355_b : _GEN_16534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16536 = 9'h164 == r_count_40_io_out ? io_r_356_b : _GEN_16535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16537 = 9'h165 == r_count_40_io_out ? io_r_357_b : _GEN_16536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16538 = 9'h166 == r_count_40_io_out ? io_r_358_b : _GEN_16537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16539 = 9'h167 == r_count_40_io_out ? io_r_359_b : _GEN_16538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16540 = 9'h168 == r_count_40_io_out ? io_r_360_b : _GEN_16539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16541 = 9'h169 == r_count_40_io_out ? io_r_361_b : _GEN_16540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16542 = 9'h16a == r_count_40_io_out ? io_r_362_b : _GEN_16541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16543 = 9'h16b == r_count_40_io_out ? io_r_363_b : _GEN_16542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16544 = 9'h16c == r_count_40_io_out ? io_r_364_b : _GEN_16543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16545 = 9'h16d == r_count_40_io_out ? io_r_365_b : _GEN_16544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16546 = 9'h16e == r_count_40_io_out ? io_r_366_b : _GEN_16545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16547 = 9'h16f == r_count_40_io_out ? io_r_367_b : _GEN_16546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16548 = 9'h170 == r_count_40_io_out ? io_r_368_b : _GEN_16547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16549 = 9'h171 == r_count_40_io_out ? io_r_369_b : _GEN_16548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16550 = 9'h172 == r_count_40_io_out ? io_r_370_b : _GEN_16549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16551 = 9'h173 == r_count_40_io_out ? io_r_371_b : _GEN_16550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16552 = 9'h174 == r_count_40_io_out ? io_r_372_b : _GEN_16551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16553 = 9'h175 == r_count_40_io_out ? io_r_373_b : _GEN_16552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16554 = 9'h176 == r_count_40_io_out ? io_r_374_b : _GEN_16553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16555 = 9'h177 == r_count_40_io_out ? io_r_375_b : _GEN_16554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16556 = 9'h178 == r_count_40_io_out ? io_r_376_b : _GEN_16555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16557 = 9'h179 == r_count_40_io_out ? io_r_377_b : _GEN_16556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16558 = 9'h17a == r_count_40_io_out ? io_r_378_b : _GEN_16557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16559 = 9'h17b == r_count_40_io_out ? io_r_379_b : _GEN_16558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16560 = 9'h17c == r_count_40_io_out ? io_r_380_b : _GEN_16559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16561 = 9'h17d == r_count_40_io_out ? io_r_381_b : _GEN_16560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16562 = 9'h17e == r_count_40_io_out ? io_r_382_b : _GEN_16561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16563 = 9'h17f == r_count_40_io_out ? io_r_383_b : _GEN_16562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16564 = 9'h180 == r_count_40_io_out ? io_r_384_b : _GEN_16563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16565 = 9'h181 == r_count_40_io_out ? io_r_385_b : _GEN_16564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16566 = 9'h182 == r_count_40_io_out ? io_r_386_b : _GEN_16565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16567 = 9'h183 == r_count_40_io_out ? io_r_387_b : _GEN_16566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16568 = 9'h184 == r_count_40_io_out ? io_r_388_b : _GEN_16567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16569 = 9'h185 == r_count_40_io_out ? io_r_389_b : _GEN_16568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16570 = 9'h186 == r_count_40_io_out ? io_r_390_b : _GEN_16569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16571 = 9'h187 == r_count_40_io_out ? io_r_391_b : _GEN_16570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16572 = 9'h188 == r_count_40_io_out ? io_r_392_b : _GEN_16571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16573 = 9'h189 == r_count_40_io_out ? io_r_393_b : _GEN_16572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16574 = 9'h18a == r_count_40_io_out ? io_r_394_b : _GEN_16573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16575 = 9'h18b == r_count_40_io_out ? io_r_395_b : _GEN_16574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16576 = 9'h18c == r_count_40_io_out ? io_r_396_b : _GEN_16575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16577 = 9'h18d == r_count_40_io_out ? io_r_397_b : _GEN_16576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16578 = 9'h18e == r_count_40_io_out ? io_r_398_b : _GEN_16577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16581 = 9'h1 == r_count_41_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16582 = 9'h2 == r_count_41_io_out ? io_r_2_b : _GEN_16581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16583 = 9'h3 == r_count_41_io_out ? io_r_3_b : _GEN_16582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16584 = 9'h4 == r_count_41_io_out ? io_r_4_b : _GEN_16583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16585 = 9'h5 == r_count_41_io_out ? io_r_5_b : _GEN_16584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16586 = 9'h6 == r_count_41_io_out ? io_r_6_b : _GEN_16585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16587 = 9'h7 == r_count_41_io_out ? io_r_7_b : _GEN_16586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16588 = 9'h8 == r_count_41_io_out ? io_r_8_b : _GEN_16587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16589 = 9'h9 == r_count_41_io_out ? io_r_9_b : _GEN_16588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16590 = 9'ha == r_count_41_io_out ? io_r_10_b : _GEN_16589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16591 = 9'hb == r_count_41_io_out ? io_r_11_b : _GEN_16590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16592 = 9'hc == r_count_41_io_out ? io_r_12_b : _GEN_16591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16593 = 9'hd == r_count_41_io_out ? io_r_13_b : _GEN_16592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16594 = 9'he == r_count_41_io_out ? io_r_14_b : _GEN_16593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16595 = 9'hf == r_count_41_io_out ? io_r_15_b : _GEN_16594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16596 = 9'h10 == r_count_41_io_out ? io_r_16_b : _GEN_16595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16597 = 9'h11 == r_count_41_io_out ? io_r_17_b : _GEN_16596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16598 = 9'h12 == r_count_41_io_out ? io_r_18_b : _GEN_16597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16599 = 9'h13 == r_count_41_io_out ? io_r_19_b : _GEN_16598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16600 = 9'h14 == r_count_41_io_out ? io_r_20_b : _GEN_16599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16601 = 9'h15 == r_count_41_io_out ? io_r_21_b : _GEN_16600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16602 = 9'h16 == r_count_41_io_out ? io_r_22_b : _GEN_16601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16603 = 9'h17 == r_count_41_io_out ? io_r_23_b : _GEN_16602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16604 = 9'h18 == r_count_41_io_out ? io_r_24_b : _GEN_16603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16605 = 9'h19 == r_count_41_io_out ? io_r_25_b : _GEN_16604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16606 = 9'h1a == r_count_41_io_out ? io_r_26_b : _GEN_16605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16607 = 9'h1b == r_count_41_io_out ? io_r_27_b : _GEN_16606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16608 = 9'h1c == r_count_41_io_out ? io_r_28_b : _GEN_16607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16609 = 9'h1d == r_count_41_io_out ? io_r_29_b : _GEN_16608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16610 = 9'h1e == r_count_41_io_out ? io_r_30_b : _GEN_16609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16611 = 9'h1f == r_count_41_io_out ? io_r_31_b : _GEN_16610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16612 = 9'h20 == r_count_41_io_out ? io_r_32_b : _GEN_16611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16613 = 9'h21 == r_count_41_io_out ? io_r_33_b : _GEN_16612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16614 = 9'h22 == r_count_41_io_out ? io_r_34_b : _GEN_16613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16615 = 9'h23 == r_count_41_io_out ? io_r_35_b : _GEN_16614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16616 = 9'h24 == r_count_41_io_out ? io_r_36_b : _GEN_16615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16617 = 9'h25 == r_count_41_io_out ? io_r_37_b : _GEN_16616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16618 = 9'h26 == r_count_41_io_out ? io_r_38_b : _GEN_16617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16619 = 9'h27 == r_count_41_io_out ? io_r_39_b : _GEN_16618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16620 = 9'h28 == r_count_41_io_out ? io_r_40_b : _GEN_16619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16621 = 9'h29 == r_count_41_io_out ? io_r_41_b : _GEN_16620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16622 = 9'h2a == r_count_41_io_out ? io_r_42_b : _GEN_16621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16623 = 9'h2b == r_count_41_io_out ? io_r_43_b : _GEN_16622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16624 = 9'h2c == r_count_41_io_out ? io_r_44_b : _GEN_16623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16625 = 9'h2d == r_count_41_io_out ? io_r_45_b : _GEN_16624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16626 = 9'h2e == r_count_41_io_out ? io_r_46_b : _GEN_16625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16627 = 9'h2f == r_count_41_io_out ? io_r_47_b : _GEN_16626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16628 = 9'h30 == r_count_41_io_out ? io_r_48_b : _GEN_16627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16629 = 9'h31 == r_count_41_io_out ? io_r_49_b : _GEN_16628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16630 = 9'h32 == r_count_41_io_out ? io_r_50_b : _GEN_16629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16631 = 9'h33 == r_count_41_io_out ? io_r_51_b : _GEN_16630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16632 = 9'h34 == r_count_41_io_out ? io_r_52_b : _GEN_16631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16633 = 9'h35 == r_count_41_io_out ? io_r_53_b : _GEN_16632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16634 = 9'h36 == r_count_41_io_out ? io_r_54_b : _GEN_16633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16635 = 9'h37 == r_count_41_io_out ? io_r_55_b : _GEN_16634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16636 = 9'h38 == r_count_41_io_out ? io_r_56_b : _GEN_16635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16637 = 9'h39 == r_count_41_io_out ? io_r_57_b : _GEN_16636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16638 = 9'h3a == r_count_41_io_out ? io_r_58_b : _GEN_16637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16639 = 9'h3b == r_count_41_io_out ? io_r_59_b : _GEN_16638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16640 = 9'h3c == r_count_41_io_out ? io_r_60_b : _GEN_16639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16641 = 9'h3d == r_count_41_io_out ? io_r_61_b : _GEN_16640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16642 = 9'h3e == r_count_41_io_out ? io_r_62_b : _GEN_16641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16643 = 9'h3f == r_count_41_io_out ? io_r_63_b : _GEN_16642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16644 = 9'h40 == r_count_41_io_out ? io_r_64_b : _GEN_16643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16645 = 9'h41 == r_count_41_io_out ? io_r_65_b : _GEN_16644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16646 = 9'h42 == r_count_41_io_out ? io_r_66_b : _GEN_16645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16647 = 9'h43 == r_count_41_io_out ? io_r_67_b : _GEN_16646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16648 = 9'h44 == r_count_41_io_out ? io_r_68_b : _GEN_16647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16649 = 9'h45 == r_count_41_io_out ? io_r_69_b : _GEN_16648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16650 = 9'h46 == r_count_41_io_out ? io_r_70_b : _GEN_16649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16651 = 9'h47 == r_count_41_io_out ? io_r_71_b : _GEN_16650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16652 = 9'h48 == r_count_41_io_out ? io_r_72_b : _GEN_16651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16653 = 9'h49 == r_count_41_io_out ? io_r_73_b : _GEN_16652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16654 = 9'h4a == r_count_41_io_out ? io_r_74_b : _GEN_16653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16655 = 9'h4b == r_count_41_io_out ? io_r_75_b : _GEN_16654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16656 = 9'h4c == r_count_41_io_out ? io_r_76_b : _GEN_16655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16657 = 9'h4d == r_count_41_io_out ? io_r_77_b : _GEN_16656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16658 = 9'h4e == r_count_41_io_out ? io_r_78_b : _GEN_16657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16659 = 9'h4f == r_count_41_io_out ? io_r_79_b : _GEN_16658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16660 = 9'h50 == r_count_41_io_out ? io_r_80_b : _GEN_16659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16661 = 9'h51 == r_count_41_io_out ? io_r_81_b : _GEN_16660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16662 = 9'h52 == r_count_41_io_out ? io_r_82_b : _GEN_16661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16663 = 9'h53 == r_count_41_io_out ? io_r_83_b : _GEN_16662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16664 = 9'h54 == r_count_41_io_out ? io_r_84_b : _GEN_16663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16665 = 9'h55 == r_count_41_io_out ? io_r_85_b : _GEN_16664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16666 = 9'h56 == r_count_41_io_out ? io_r_86_b : _GEN_16665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16667 = 9'h57 == r_count_41_io_out ? io_r_87_b : _GEN_16666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16668 = 9'h58 == r_count_41_io_out ? io_r_88_b : _GEN_16667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16669 = 9'h59 == r_count_41_io_out ? io_r_89_b : _GEN_16668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16670 = 9'h5a == r_count_41_io_out ? io_r_90_b : _GEN_16669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16671 = 9'h5b == r_count_41_io_out ? io_r_91_b : _GEN_16670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16672 = 9'h5c == r_count_41_io_out ? io_r_92_b : _GEN_16671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16673 = 9'h5d == r_count_41_io_out ? io_r_93_b : _GEN_16672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16674 = 9'h5e == r_count_41_io_out ? io_r_94_b : _GEN_16673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16675 = 9'h5f == r_count_41_io_out ? io_r_95_b : _GEN_16674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16676 = 9'h60 == r_count_41_io_out ? io_r_96_b : _GEN_16675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16677 = 9'h61 == r_count_41_io_out ? io_r_97_b : _GEN_16676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16678 = 9'h62 == r_count_41_io_out ? io_r_98_b : _GEN_16677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16679 = 9'h63 == r_count_41_io_out ? io_r_99_b : _GEN_16678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16680 = 9'h64 == r_count_41_io_out ? io_r_100_b : _GEN_16679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16681 = 9'h65 == r_count_41_io_out ? io_r_101_b : _GEN_16680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16682 = 9'h66 == r_count_41_io_out ? io_r_102_b : _GEN_16681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16683 = 9'h67 == r_count_41_io_out ? io_r_103_b : _GEN_16682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16684 = 9'h68 == r_count_41_io_out ? io_r_104_b : _GEN_16683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16685 = 9'h69 == r_count_41_io_out ? io_r_105_b : _GEN_16684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16686 = 9'h6a == r_count_41_io_out ? io_r_106_b : _GEN_16685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16687 = 9'h6b == r_count_41_io_out ? io_r_107_b : _GEN_16686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16688 = 9'h6c == r_count_41_io_out ? io_r_108_b : _GEN_16687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16689 = 9'h6d == r_count_41_io_out ? io_r_109_b : _GEN_16688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16690 = 9'h6e == r_count_41_io_out ? io_r_110_b : _GEN_16689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16691 = 9'h6f == r_count_41_io_out ? io_r_111_b : _GEN_16690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16692 = 9'h70 == r_count_41_io_out ? io_r_112_b : _GEN_16691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16693 = 9'h71 == r_count_41_io_out ? io_r_113_b : _GEN_16692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16694 = 9'h72 == r_count_41_io_out ? io_r_114_b : _GEN_16693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16695 = 9'h73 == r_count_41_io_out ? io_r_115_b : _GEN_16694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16696 = 9'h74 == r_count_41_io_out ? io_r_116_b : _GEN_16695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16697 = 9'h75 == r_count_41_io_out ? io_r_117_b : _GEN_16696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16698 = 9'h76 == r_count_41_io_out ? io_r_118_b : _GEN_16697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16699 = 9'h77 == r_count_41_io_out ? io_r_119_b : _GEN_16698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16700 = 9'h78 == r_count_41_io_out ? io_r_120_b : _GEN_16699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16701 = 9'h79 == r_count_41_io_out ? io_r_121_b : _GEN_16700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16702 = 9'h7a == r_count_41_io_out ? io_r_122_b : _GEN_16701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16703 = 9'h7b == r_count_41_io_out ? io_r_123_b : _GEN_16702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16704 = 9'h7c == r_count_41_io_out ? io_r_124_b : _GEN_16703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16705 = 9'h7d == r_count_41_io_out ? io_r_125_b : _GEN_16704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16706 = 9'h7e == r_count_41_io_out ? io_r_126_b : _GEN_16705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16707 = 9'h7f == r_count_41_io_out ? io_r_127_b : _GEN_16706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16708 = 9'h80 == r_count_41_io_out ? io_r_128_b : _GEN_16707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16709 = 9'h81 == r_count_41_io_out ? io_r_129_b : _GEN_16708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16710 = 9'h82 == r_count_41_io_out ? io_r_130_b : _GEN_16709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16711 = 9'h83 == r_count_41_io_out ? io_r_131_b : _GEN_16710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16712 = 9'h84 == r_count_41_io_out ? io_r_132_b : _GEN_16711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16713 = 9'h85 == r_count_41_io_out ? io_r_133_b : _GEN_16712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16714 = 9'h86 == r_count_41_io_out ? io_r_134_b : _GEN_16713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16715 = 9'h87 == r_count_41_io_out ? io_r_135_b : _GEN_16714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16716 = 9'h88 == r_count_41_io_out ? io_r_136_b : _GEN_16715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16717 = 9'h89 == r_count_41_io_out ? io_r_137_b : _GEN_16716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16718 = 9'h8a == r_count_41_io_out ? io_r_138_b : _GEN_16717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16719 = 9'h8b == r_count_41_io_out ? io_r_139_b : _GEN_16718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16720 = 9'h8c == r_count_41_io_out ? io_r_140_b : _GEN_16719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16721 = 9'h8d == r_count_41_io_out ? io_r_141_b : _GEN_16720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16722 = 9'h8e == r_count_41_io_out ? io_r_142_b : _GEN_16721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16723 = 9'h8f == r_count_41_io_out ? io_r_143_b : _GEN_16722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16724 = 9'h90 == r_count_41_io_out ? io_r_144_b : _GEN_16723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16725 = 9'h91 == r_count_41_io_out ? io_r_145_b : _GEN_16724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16726 = 9'h92 == r_count_41_io_out ? io_r_146_b : _GEN_16725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16727 = 9'h93 == r_count_41_io_out ? io_r_147_b : _GEN_16726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16728 = 9'h94 == r_count_41_io_out ? io_r_148_b : _GEN_16727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16729 = 9'h95 == r_count_41_io_out ? io_r_149_b : _GEN_16728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16730 = 9'h96 == r_count_41_io_out ? io_r_150_b : _GEN_16729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16731 = 9'h97 == r_count_41_io_out ? io_r_151_b : _GEN_16730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16732 = 9'h98 == r_count_41_io_out ? io_r_152_b : _GEN_16731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16733 = 9'h99 == r_count_41_io_out ? io_r_153_b : _GEN_16732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16734 = 9'h9a == r_count_41_io_out ? io_r_154_b : _GEN_16733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16735 = 9'h9b == r_count_41_io_out ? io_r_155_b : _GEN_16734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16736 = 9'h9c == r_count_41_io_out ? io_r_156_b : _GEN_16735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16737 = 9'h9d == r_count_41_io_out ? io_r_157_b : _GEN_16736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16738 = 9'h9e == r_count_41_io_out ? io_r_158_b : _GEN_16737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16739 = 9'h9f == r_count_41_io_out ? io_r_159_b : _GEN_16738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16740 = 9'ha0 == r_count_41_io_out ? io_r_160_b : _GEN_16739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16741 = 9'ha1 == r_count_41_io_out ? io_r_161_b : _GEN_16740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16742 = 9'ha2 == r_count_41_io_out ? io_r_162_b : _GEN_16741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16743 = 9'ha3 == r_count_41_io_out ? io_r_163_b : _GEN_16742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16744 = 9'ha4 == r_count_41_io_out ? io_r_164_b : _GEN_16743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16745 = 9'ha5 == r_count_41_io_out ? io_r_165_b : _GEN_16744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16746 = 9'ha6 == r_count_41_io_out ? io_r_166_b : _GEN_16745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16747 = 9'ha7 == r_count_41_io_out ? io_r_167_b : _GEN_16746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16748 = 9'ha8 == r_count_41_io_out ? io_r_168_b : _GEN_16747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16749 = 9'ha9 == r_count_41_io_out ? io_r_169_b : _GEN_16748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16750 = 9'haa == r_count_41_io_out ? io_r_170_b : _GEN_16749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16751 = 9'hab == r_count_41_io_out ? io_r_171_b : _GEN_16750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16752 = 9'hac == r_count_41_io_out ? io_r_172_b : _GEN_16751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16753 = 9'had == r_count_41_io_out ? io_r_173_b : _GEN_16752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16754 = 9'hae == r_count_41_io_out ? io_r_174_b : _GEN_16753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16755 = 9'haf == r_count_41_io_out ? io_r_175_b : _GEN_16754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16756 = 9'hb0 == r_count_41_io_out ? io_r_176_b : _GEN_16755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16757 = 9'hb1 == r_count_41_io_out ? io_r_177_b : _GEN_16756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16758 = 9'hb2 == r_count_41_io_out ? io_r_178_b : _GEN_16757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16759 = 9'hb3 == r_count_41_io_out ? io_r_179_b : _GEN_16758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16760 = 9'hb4 == r_count_41_io_out ? io_r_180_b : _GEN_16759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16761 = 9'hb5 == r_count_41_io_out ? io_r_181_b : _GEN_16760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16762 = 9'hb6 == r_count_41_io_out ? io_r_182_b : _GEN_16761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16763 = 9'hb7 == r_count_41_io_out ? io_r_183_b : _GEN_16762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16764 = 9'hb8 == r_count_41_io_out ? io_r_184_b : _GEN_16763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16765 = 9'hb9 == r_count_41_io_out ? io_r_185_b : _GEN_16764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16766 = 9'hba == r_count_41_io_out ? io_r_186_b : _GEN_16765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16767 = 9'hbb == r_count_41_io_out ? io_r_187_b : _GEN_16766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16768 = 9'hbc == r_count_41_io_out ? io_r_188_b : _GEN_16767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16769 = 9'hbd == r_count_41_io_out ? io_r_189_b : _GEN_16768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16770 = 9'hbe == r_count_41_io_out ? io_r_190_b : _GEN_16769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16771 = 9'hbf == r_count_41_io_out ? io_r_191_b : _GEN_16770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16772 = 9'hc0 == r_count_41_io_out ? io_r_192_b : _GEN_16771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16773 = 9'hc1 == r_count_41_io_out ? io_r_193_b : _GEN_16772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16774 = 9'hc2 == r_count_41_io_out ? io_r_194_b : _GEN_16773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16775 = 9'hc3 == r_count_41_io_out ? io_r_195_b : _GEN_16774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16776 = 9'hc4 == r_count_41_io_out ? io_r_196_b : _GEN_16775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16777 = 9'hc5 == r_count_41_io_out ? io_r_197_b : _GEN_16776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16778 = 9'hc6 == r_count_41_io_out ? io_r_198_b : _GEN_16777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16779 = 9'hc7 == r_count_41_io_out ? io_r_199_b : _GEN_16778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16780 = 9'hc8 == r_count_41_io_out ? io_r_200_b : _GEN_16779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16781 = 9'hc9 == r_count_41_io_out ? io_r_201_b : _GEN_16780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16782 = 9'hca == r_count_41_io_out ? io_r_202_b : _GEN_16781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16783 = 9'hcb == r_count_41_io_out ? io_r_203_b : _GEN_16782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16784 = 9'hcc == r_count_41_io_out ? io_r_204_b : _GEN_16783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16785 = 9'hcd == r_count_41_io_out ? io_r_205_b : _GEN_16784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16786 = 9'hce == r_count_41_io_out ? io_r_206_b : _GEN_16785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16787 = 9'hcf == r_count_41_io_out ? io_r_207_b : _GEN_16786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16788 = 9'hd0 == r_count_41_io_out ? io_r_208_b : _GEN_16787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16789 = 9'hd1 == r_count_41_io_out ? io_r_209_b : _GEN_16788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16790 = 9'hd2 == r_count_41_io_out ? io_r_210_b : _GEN_16789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16791 = 9'hd3 == r_count_41_io_out ? io_r_211_b : _GEN_16790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16792 = 9'hd4 == r_count_41_io_out ? io_r_212_b : _GEN_16791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16793 = 9'hd5 == r_count_41_io_out ? io_r_213_b : _GEN_16792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16794 = 9'hd6 == r_count_41_io_out ? io_r_214_b : _GEN_16793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16795 = 9'hd7 == r_count_41_io_out ? io_r_215_b : _GEN_16794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16796 = 9'hd8 == r_count_41_io_out ? io_r_216_b : _GEN_16795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16797 = 9'hd9 == r_count_41_io_out ? io_r_217_b : _GEN_16796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16798 = 9'hda == r_count_41_io_out ? io_r_218_b : _GEN_16797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16799 = 9'hdb == r_count_41_io_out ? io_r_219_b : _GEN_16798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16800 = 9'hdc == r_count_41_io_out ? io_r_220_b : _GEN_16799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16801 = 9'hdd == r_count_41_io_out ? io_r_221_b : _GEN_16800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16802 = 9'hde == r_count_41_io_out ? io_r_222_b : _GEN_16801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16803 = 9'hdf == r_count_41_io_out ? io_r_223_b : _GEN_16802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16804 = 9'he0 == r_count_41_io_out ? io_r_224_b : _GEN_16803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16805 = 9'he1 == r_count_41_io_out ? io_r_225_b : _GEN_16804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16806 = 9'he2 == r_count_41_io_out ? io_r_226_b : _GEN_16805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16807 = 9'he3 == r_count_41_io_out ? io_r_227_b : _GEN_16806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16808 = 9'he4 == r_count_41_io_out ? io_r_228_b : _GEN_16807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16809 = 9'he5 == r_count_41_io_out ? io_r_229_b : _GEN_16808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16810 = 9'he6 == r_count_41_io_out ? io_r_230_b : _GEN_16809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16811 = 9'he7 == r_count_41_io_out ? io_r_231_b : _GEN_16810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16812 = 9'he8 == r_count_41_io_out ? io_r_232_b : _GEN_16811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16813 = 9'he9 == r_count_41_io_out ? io_r_233_b : _GEN_16812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16814 = 9'hea == r_count_41_io_out ? io_r_234_b : _GEN_16813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16815 = 9'heb == r_count_41_io_out ? io_r_235_b : _GEN_16814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16816 = 9'hec == r_count_41_io_out ? io_r_236_b : _GEN_16815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16817 = 9'hed == r_count_41_io_out ? io_r_237_b : _GEN_16816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16818 = 9'hee == r_count_41_io_out ? io_r_238_b : _GEN_16817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16819 = 9'hef == r_count_41_io_out ? io_r_239_b : _GEN_16818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16820 = 9'hf0 == r_count_41_io_out ? io_r_240_b : _GEN_16819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16821 = 9'hf1 == r_count_41_io_out ? io_r_241_b : _GEN_16820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16822 = 9'hf2 == r_count_41_io_out ? io_r_242_b : _GEN_16821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16823 = 9'hf3 == r_count_41_io_out ? io_r_243_b : _GEN_16822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16824 = 9'hf4 == r_count_41_io_out ? io_r_244_b : _GEN_16823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16825 = 9'hf5 == r_count_41_io_out ? io_r_245_b : _GEN_16824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16826 = 9'hf6 == r_count_41_io_out ? io_r_246_b : _GEN_16825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16827 = 9'hf7 == r_count_41_io_out ? io_r_247_b : _GEN_16826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16828 = 9'hf8 == r_count_41_io_out ? io_r_248_b : _GEN_16827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16829 = 9'hf9 == r_count_41_io_out ? io_r_249_b : _GEN_16828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16830 = 9'hfa == r_count_41_io_out ? io_r_250_b : _GEN_16829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16831 = 9'hfb == r_count_41_io_out ? io_r_251_b : _GEN_16830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16832 = 9'hfc == r_count_41_io_out ? io_r_252_b : _GEN_16831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16833 = 9'hfd == r_count_41_io_out ? io_r_253_b : _GEN_16832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16834 = 9'hfe == r_count_41_io_out ? io_r_254_b : _GEN_16833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16835 = 9'hff == r_count_41_io_out ? io_r_255_b : _GEN_16834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16836 = 9'h100 == r_count_41_io_out ? io_r_256_b : _GEN_16835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16837 = 9'h101 == r_count_41_io_out ? io_r_257_b : _GEN_16836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16838 = 9'h102 == r_count_41_io_out ? io_r_258_b : _GEN_16837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16839 = 9'h103 == r_count_41_io_out ? io_r_259_b : _GEN_16838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16840 = 9'h104 == r_count_41_io_out ? io_r_260_b : _GEN_16839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16841 = 9'h105 == r_count_41_io_out ? io_r_261_b : _GEN_16840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16842 = 9'h106 == r_count_41_io_out ? io_r_262_b : _GEN_16841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16843 = 9'h107 == r_count_41_io_out ? io_r_263_b : _GEN_16842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16844 = 9'h108 == r_count_41_io_out ? io_r_264_b : _GEN_16843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16845 = 9'h109 == r_count_41_io_out ? io_r_265_b : _GEN_16844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16846 = 9'h10a == r_count_41_io_out ? io_r_266_b : _GEN_16845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16847 = 9'h10b == r_count_41_io_out ? io_r_267_b : _GEN_16846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16848 = 9'h10c == r_count_41_io_out ? io_r_268_b : _GEN_16847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16849 = 9'h10d == r_count_41_io_out ? io_r_269_b : _GEN_16848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16850 = 9'h10e == r_count_41_io_out ? io_r_270_b : _GEN_16849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16851 = 9'h10f == r_count_41_io_out ? io_r_271_b : _GEN_16850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16852 = 9'h110 == r_count_41_io_out ? io_r_272_b : _GEN_16851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16853 = 9'h111 == r_count_41_io_out ? io_r_273_b : _GEN_16852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16854 = 9'h112 == r_count_41_io_out ? io_r_274_b : _GEN_16853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16855 = 9'h113 == r_count_41_io_out ? io_r_275_b : _GEN_16854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16856 = 9'h114 == r_count_41_io_out ? io_r_276_b : _GEN_16855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16857 = 9'h115 == r_count_41_io_out ? io_r_277_b : _GEN_16856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16858 = 9'h116 == r_count_41_io_out ? io_r_278_b : _GEN_16857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16859 = 9'h117 == r_count_41_io_out ? io_r_279_b : _GEN_16858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16860 = 9'h118 == r_count_41_io_out ? io_r_280_b : _GEN_16859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16861 = 9'h119 == r_count_41_io_out ? io_r_281_b : _GEN_16860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16862 = 9'h11a == r_count_41_io_out ? io_r_282_b : _GEN_16861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16863 = 9'h11b == r_count_41_io_out ? io_r_283_b : _GEN_16862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16864 = 9'h11c == r_count_41_io_out ? io_r_284_b : _GEN_16863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16865 = 9'h11d == r_count_41_io_out ? io_r_285_b : _GEN_16864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16866 = 9'h11e == r_count_41_io_out ? io_r_286_b : _GEN_16865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16867 = 9'h11f == r_count_41_io_out ? io_r_287_b : _GEN_16866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16868 = 9'h120 == r_count_41_io_out ? io_r_288_b : _GEN_16867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16869 = 9'h121 == r_count_41_io_out ? io_r_289_b : _GEN_16868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16870 = 9'h122 == r_count_41_io_out ? io_r_290_b : _GEN_16869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16871 = 9'h123 == r_count_41_io_out ? io_r_291_b : _GEN_16870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16872 = 9'h124 == r_count_41_io_out ? io_r_292_b : _GEN_16871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16873 = 9'h125 == r_count_41_io_out ? io_r_293_b : _GEN_16872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16874 = 9'h126 == r_count_41_io_out ? io_r_294_b : _GEN_16873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16875 = 9'h127 == r_count_41_io_out ? io_r_295_b : _GEN_16874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16876 = 9'h128 == r_count_41_io_out ? io_r_296_b : _GEN_16875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16877 = 9'h129 == r_count_41_io_out ? io_r_297_b : _GEN_16876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16878 = 9'h12a == r_count_41_io_out ? io_r_298_b : _GEN_16877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16879 = 9'h12b == r_count_41_io_out ? io_r_299_b : _GEN_16878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16880 = 9'h12c == r_count_41_io_out ? io_r_300_b : _GEN_16879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16881 = 9'h12d == r_count_41_io_out ? io_r_301_b : _GEN_16880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16882 = 9'h12e == r_count_41_io_out ? io_r_302_b : _GEN_16881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16883 = 9'h12f == r_count_41_io_out ? io_r_303_b : _GEN_16882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16884 = 9'h130 == r_count_41_io_out ? io_r_304_b : _GEN_16883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16885 = 9'h131 == r_count_41_io_out ? io_r_305_b : _GEN_16884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16886 = 9'h132 == r_count_41_io_out ? io_r_306_b : _GEN_16885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16887 = 9'h133 == r_count_41_io_out ? io_r_307_b : _GEN_16886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16888 = 9'h134 == r_count_41_io_out ? io_r_308_b : _GEN_16887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16889 = 9'h135 == r_count_41_io_out ? io_r_309_b : _GEN_16888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16890 = 9'h136 == r_count_41_io_out ? io_r_310_b : _GEN_16889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16891 = 9'h137 == r_count_41_io_out ? io_r_311_b : _GEN_16890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16892 = 9'h138 == r_count_41_io_out ? io_r_312_b : _GEN_16891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16893 = 9'h139 == r_count_41_io_out ? io_r_313_b : _GEN_16892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16894 = 9'h13a == r_count_41_io_out ? io_r_314_b : _GEN_16893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16895 = 9'h13b == r_count_41_io_out ? io_r_315_b : _GEN_16894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16896 = 9'h13c == r_count_41_io_out ? io_r_316_b : _GEN_16895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16897 = 9'h13d == r_count_41_io_out ? io_r_317_b : _GEN_16896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16898 = 9'h13e == r_count_41_io_out ? io_r_318_b : _GEN_16897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16899 = 9'h13f == r_count_41_io_out ? io_r_319_b : _GEN_16898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16900 = 9'h140 == r_count_41_io_out ? io_r_320_b : _GEN_16899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16901 = 9'h141 == r_count_41_io_out ? io_r_321_b : _GEN_16900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16902 = 9'h142 == r_count_41_io_out ? io_r_322_b : _GEN_16901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16903 = 9'h143 == r_count_41_io_out ? io_r_323_b : _GEN_16902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16904 = 9'h144 == r_count_41_io_out ? io_r_324_b : _GEN_16903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16905 = 9'h145 == r_count_41_io_out ? io_r_325_b : _GEN_16904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16906 = 9'h146 == r_count_41_io_out ? io_r_326_b : _GEN_16905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16907 = 9'h147 == r_count_41_io_out ? io_r_327_b : _GEN_16906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16908 = 9'h148 == r_count_41_io_out ? io_r_328_b : _GEN_16907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16909 = 9'h149 == r_count_41_io_out ? io_r_329_b : _GEN_16908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16910 = 9'h14a == r_count_41_io_out ? io_r_330_b : _GEN_16909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16911 = 9'h14b == r_count_41_io_out ? io_r_331_b : _GEN_16910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16912 = 9'h14c == r_count_41_io_out ? io_r_332_b : _GEN_16911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16913 = 9'h14d == r_count_41_io_out ? io_r_333_b : _GEN_16912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16914 = 9'h14e == r_count_41_io_out ? io_r_334_b : _GEN_16913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16915 = 9'h14f == r_count_41_io_out ? io_r_335_b : _GEN_16914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16916 = 9'h150 == r_count_41_io_out ? io_r_336_b : _GEN_16915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16917 = 9'h151 == r_count_41_io_out ? io_r_337_b : _GEN_16916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16918 = 9'h152 == r_count_41_io_out ? io_r_338_b : _GEN_16917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16919 = 9'h153 == r_count_41_io_out ? io_r_339_b : _GEN_16918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16920 = 9'h154 == r_count_41_io_out ? io_r_340_b : _GEN_16919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16921 = 9'h155 == r_count_41_io_out ? io_r_341_b : _GEN_16920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16922 = 9'h156 == r_count_41_io_out ? io_r_342_b : _GEN_16921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16923 = 9'h157 == r_count_41_io_out ? io_r_343_b : _GEN_16922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16924 = 9'h158 == r_count_41_io_out ? io_r_344_b : _GEN_16923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16925 = 9'h159 == r_count_41_io_out ? io_r_345_b : _GEN_16924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16926 = 9'h15a == r_count_41_io_out ? io_r_346_b : _GEN_16925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16927 = 9'h15b == r_count_41_io_out ? io_r_347_b : _GEN_16926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16928 = 9'h15c == r_count_41_io_out ? io_r_348_b : _GEN_16927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16929 = 9'h15d == r_count_41_io_out ? io_r_349_b : _GEN_16928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16930 = 9'h15e == r_count_41_io_out ? io_r_350_b : _GEN_16929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16931 = 9'h15f == r_count_41_io_out ? io_r_351_b : _GEN_16930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16932 = 9'h160 == r_count_41_io_out ? io_r_352_b : _GEN_16931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16933 = 9'h161 == r_count_41_io_out ? io_r_353_b : _GEN_16932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16934 = 9'h162 == r_count_41_io_out ? io_r_354_b : _GEN_16933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16935 = 9'h163 == r_count_41_io_out ? io_r_355_b : _GEN_16934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16936 = 9'h164 == r_count_41_io_out ? io_r_356_b : _GEN_16935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16937 = 9'h165 == r_count_41_io_out ? io_r_357_b : _GEN_16936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16938 = 9'h166 == r_count_41_io_out ? io_r_358_b : _GEN_16937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16939 = 9'h167 == r_count_41_io_out ? io_r_359_b : _GEN_16938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16940 = 9'h168 == r_count_41_io_out ? io_r_360_b : _GEN_16939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16941 = 9'h169 == r_count_41_io_out ? io_r_361_b : _GEN_16940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16942 = 9'h16a == r_count_41_io_out ? io_r_362_b : _GEN_16941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16943 = 9'h16b == r_count_41_io_out ? io_r_363_b : _GEN_16942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16944 = 9'h16c == r_count_41_io_out ? io_r_364_b : _GEN_16943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16945 = 9'h16d == r_count_41_io_out ? io_r_365_b : _GEN_16944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16946 = 9'h16e == r_count_41_io_out ? io_r_366_b : _GEN_16945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16947 = 9'h16f == r_count_41_io_out ? io_r_367_b : _GEN_16946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16948 = 9'h170 == r_count_41_io_out ? io_r_368_b : _GEN_16947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16949 = 9'h171 == r_count_41_io_out ? io_r_369_b : _GEN_16948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16950 = 9'h172 == r_count_41_io_out ? io_r_370_b : _GEN_16949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16951 = 9'h173 == r_count_41_io_out ? io_r_371_b : _GEN_16950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16952 = 9'h174 == r_count_41_io_out ? io_r_372_b : _GEN_16951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16953 = 9'h175 == r_count_41_io_out ? io_r_373_b : _GEN_16952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16954 = 9'h176 == r_count_41_io_out ? io_r_374_b : _GEN_16953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16955 = 9'h177 == r_count_41_io_out ? io_r_375_b : _GEN_16954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16956 = 9'h178 == r_count_41_io_out ? io_r_376_b : _GEN_16955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16957 = 9'h179 == r_count_41_io_out ? io_r_377_b : _GEN_16956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16958 = 9'h17a == r_count_41_io_out ? io_r_378_b : _GEN_16957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16959 = 9'h17b == r_count_41_io_out ? io_r_379_b : _GEN_16958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16960 = 9'h17c == r_count_41_io_out ? io_r_380_b : _GEN_16959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16961 = 9'h17d == r_count_41_io_out ? io_r_381_b : _GEN_16960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16962 = 9'h17e == r_count_41_io_out ? io_r_382_b : _GEN_16961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16963 = 9'h17f == r_count_41_io_out ? io_r_383_b : _GEN_16962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16964 = 9'h180 == r_count_41_io_out ? io_r_384_b : _GEN_16963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16965 = 9'h181 == r_count_41_io_out ? io_r_385_b : _GEN_16964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16966 = 9'h182 == r_count_41_io_out ? io_r_386_b : _GEN_16965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16967 = 9'h183 == r_count_41_io_out ? io_r_387_b : _GEN_16966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16968 = 9'h184 == r_count_41_io_out ? io_r_388_b : _GEN_16967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16969 = 9'h185 == r_count_41_io_out ? io_r_389_b : _GEN_16968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16970 = 9'h186 == r_count_41_io_out ? io_r_390_b : _GEN_16969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16971 = 9'h187 == r_count_41_io_out ? io_r_391_b : _GEN_16970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16972 = 9'h188 == r_count_41_io_out ? io_r_392_b : _GEN_16971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16973 = 9'h189 == r_count_41_io_out ? io_r_393_b : _GEN_16972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16974 = 9'h18a == r_count_41_io_out ? io_r_394_b : _GEN_16973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16975 = 9'h18b == r_count_41_io_out ? io_r_395_b : _GEN_16974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16976 = 9'h18c == r_count_41_io_out ? io_r_396_b : _GEN_16975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16977 = 9'h18d == r_count_41_io_out ? io_r_397_b : _GEN_16976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16978 = 9'h18e == r_count_41_io_out ? io_r_398_b : _GEN_16977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16981 = 9'h1 == r_count_42_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16982 = 9'h2 == r_count_42_io_out ? io_r_2_b : _GEN_16981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16983 = 9'h3 == r_count_42_io_out ? io_r_3_b : _GEN_16982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16984 = 9'h4 == r_count_42_io_out ? io_r_4_b : _GEN_16983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16985 = 9'h5 == r_count_42_io_out ? io_r_5_b : _GEN_16984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16986 = 9'h6 == r_count_42_io_out ? io_r_6_b : _GEN_16985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16987 = 9'h7 == r_count_42_io_out ? io_r_7_b : _GEN_16986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16988 = 9'h8 == r_count_42_io_out ? io_r_8_b : _GEN_16987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16989 = 9'h9 == r_count_42_io_out ? io_r_9_b : _GEN_16988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16990 = 9'ha == r_count_42_io_out ? io_r_10_b : _GEN_16989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16991 = 9'hb == r_count_42_io_out ? io_r_11_b : _GEN_16990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16992 = 9'hc == r_count_42_io_out ? io_r_12_b : _GEN_16991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16993 = 9'hd == r_count_42_io_out ? io_r_13_b : _GEN_16992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16994 = 9'he == r_count_42_io_out ? io_r_14_b : _GEN_16993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16995 = 9'hf == r_count_42_io_out ? io_r_15_b : _GEN_16994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16996 = 9'h10 == r_count_42_io_out ? io_r_16_b : _GEN_16995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16997 = 9'h11 == r_count_42_io_out ? io_r_17_b : _GEN_16996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16998 = 9'h12 == r_count_42_io_out ? io_r_18_b : _GEN_16997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16999 = 9'h13 == r_count_42_io_out ? io_r_19_b : _GEN_16998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17000 = 9'h14 == r_count_42_io_out ? io_r_20_b : _GEN_16999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17001 = 9'h15 == r_count_42_io_out ? io_r_21_b : _GEN_17000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17002 = 9'h16 == r_count_42_io_out ? io_r_22_b : _GEN_17001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17003 = 9'h17 == r_count_42_io_out ? io_r_23_b : _GEN_17002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17004 = 9'h18 == r_count_42_io_out ? io_r_24_b : _GEN_17003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17005 = 9'h19 == r_count_42_io_out ? io_r_25_b : _GEN_17004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17006 = 9'h1a == r_count_42_io_out ? io_r_26_b : _GEN_17005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17007 = 9'h1b == r_count_42_io_out ? io_r_27_b : _GEN_17006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17008 = 9'h1c == r_count_42_io_out ? io_r_28_b : _GEN_17007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17009 = 9'h1d == r_count_42_io_out ? io_r_29_b : _GEN_17008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17010 = 9'h1e == r_count_42_io_out ? io_r_30_b : _GEN_17009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17011 = 9'h1f == r_count_42_io_out ? io_r_31_b : _GEN_17010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17012 = 9'h20 == r_count_42_io_out ? io_r_32_b : _GEN_17011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17013 = 9'h21 == r_count_42_io_out ? io_r_33_b : _GEN_17012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17014 = 9'h22 == r_count_42_io_out ? io_r_34_b : _GEN_17013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17015 = 9'h23 == r_count_42_io_out ? io_r_35_b : _GEN_17014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17016 = 9'h24 == r_count_42_io_out ? io_r_36_b : _GEN_17015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17017 = 9'h25 == r_count_42_io_out ? io_r_37_b : _GEN_17016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17018 = 9'h26 == r_count_42_io_out ? io_r_38_b : _GEN_17017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17019 = 9'h27 == r_count_42_io_out ? io_r_39_b : _GEN_17018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17020 = 9'h28 == r_count_42_io_out ? io_r_40_b : _GEN_17019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17021 = 9'h29 == r_count_42_io_out ? io_r_41_b : _GEN_17020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17022 = 9'h2a == r_count_42_io_out ? io_r_42_b : _GEN_17021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17023 = 9'h2b == r_count_42_io_out ? io_r_43_b : _GEN_17022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17024 = 9'h2c == r_count_42_io_out ? io_r_44_b : _GEN_17023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17025 = 9'h2d == r_count_42_io_out ? io_r_45_b : _GEN_17024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17026 = 9'h2e == r_count_42_io_out ? io_r_46_b : _GEN_17025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17027 = 9'h2f == r_count_42_io_out ? io_r_47_b : _GEN_17026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17028 = 9'h30 == r_count_42_io_out ? io_r_48_b : _GEN_17027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17029 = 9'h31 == r_count_42_io_out ? io_r_49_b : _GEN_17028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17030 = 9'h32 == r_count_42_io_out ? io_r_50_b : _GEN_17029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17031 = 9'h33 == r_count_42_io_out ? io_r_51_b : _GEN_17030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17032 = 9'h34 == r_count_42_io_out ? io_r_52_b : _GEN_17031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17033 = 9'h35 == r_count_42_io_out ? io_r_53_b : _GEN_17032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17034 = 9'h36 == r_count_42_io_out ? io_r_54_b : _GEN_17033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17035 = 9'h37 == r_count_42_io_out ? io_r_55_b : _GEN_17034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17036 = 9'h38 == r_count_42_io_out ? io_r_56_b : _GEN_17035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17037 = 9'h39 == r_count_42_io_out ? io_r_57_b : _GEN_17036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17038 = 9'h3a == r_count_42_io_out ? io_r_58_b : _GEN_17037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17039 = 9'h3b == r_count_42_io_out ? io_r_59_b : _GEN_17038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17040 = 9'h3c == r_count_42_io_out ? io_r_60_b : _GEN_17039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17041 = 9'h3d == r_count_42_io_out ? io_r_61_b : _GEN_17040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17042 = 9'h3e == r_count_42_io_out ? io_r_62_b : _GEN_17041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17043 = 9'h3f == r_count_42_io_out ? io_r_63_b : _GEN_17042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17044 = 9'h40 == r_count_42_io_out ? io_r_64_b : _GEN_17043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17045 = 9'h41 == r_count_42_io_out ? io_r_65_b : _GEN_17044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17046 = 9'h42 == r_count_42_io_out ? io_r_66_b : _GEN_17045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17047 = 9'h43 == r_count_42_io_out ? io_r_67_b : _GEN_17046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17048 = 9'h44 == r_count_42_io_out ? io_r_68_b : _GEN_17047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17049 = 9'h45 == r_count_42_io_out ? io_r_69_b : _GEN_17048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17050 = 9'h46 == r_count_42_io_out ? io_r_70_b : _GEN_17049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17051 = 9'h47 == r_count_42_io_out ? io_r_71_b : _GEN_17050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17052 = 9'h48 == r_count_42_io_out ? io_r_72_b : _GEN_17051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17053 = 9'h49 == r_count_42_io_out ? io_r_73_b : _GEN_17052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17054 = 9'h4a == r_count_42_io_out ? io_r_74_b : _GEN_17053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17055 = 9'h4b == r_count_42_io_out ? io_r_75_b : _GEN_17054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17056 = 9'h4c == r_count_42_io_out ? io_r_76_b : _GEN_17055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17057 = 9'h4d == r_count_42_io_out ? io_r_77_b : _GEN_17056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17058 = 9'h4e == r_count_42_io_out ? io_r_78_b : _GEN_17057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17059 = 9'h4f == r_count_42_io_out ? io_r_79_b : _GEN_17058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17060 = 9'h50 == r_count_42_io_out ? io_r_80_b : _GEN_17059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17061 = 9'h51 == r_count_42_io_out ? io_r_81_b : _GEN_17060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17062 = 9'h52 == r_count_42_io_out ? io_r_82_b : _GEN_17061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17063 = 9'h53 == r_count_42_io_out ? io_r_83_b : _GEN_17062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17064 = 9'h54 == r_count_42_io_out ? io_r_84_b : _GEN_17063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17065 = 9'h55 == r_count_42_io_out ? io_r_85_b : _GEN_17064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17066 = 9'h56 == r_count_42_io_out ? io_r_86_b : _GEN_17065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17067 = 9'h57 == r_count_42_io_out ? io_r_87_b : _GEN_17066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17068 = 9'h58 == r_count_42_io_out ? io_r_88_b : _GEN_17067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17069 = 9'h59 == r_count_42_io_out ? io_r_89_b : _GEN_17068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17070 = 9'h5a == r_count_42_io_out ? io_r_90_b : _GEN_17069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17071 = 9'h5b == r_count_42_io_out ? io_r_91_b : _GEN_17070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17072 = 9'h5c == r_count_42_io_out ? io_r_92_b : _GEN_17071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17073 = 9'h5d == r_count_42_io_out ? io_r_93_b : _GEN_17072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17074 = 9'h5e == r_count_42_io_out ? io_r_94_b : _GEN_17073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17075 = 9'h5f == r_count_42_io_out ? io_r_95_b : _GEN_17074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17076 = 9'h60 == r_count_42_io_out ? io_r_96_b : _GEN_17075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17077 = 9'h61 == r_count_42_io_out ? io_r_97_b : _GEN_17076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17078 = 9'h62 == r_count_42_io_out ? io_r_98_b : _GEN_17077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17079 = 9'h63 == r_count_42_io_out ? io_r_99_b : _GEN_17078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17080 = 9'h64 == r_count_42_io_out ? io_r_100_b : _GEN_17079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17081 = 9'h65 == r_count_42_io_out ? io_r_101_b : _GEN_17080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17082 = 9'h66 == r_count_42_io_out ? io_r_102_b : _GEN_17081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17083 = 9'h67 == r_count_42_io_out ? io_r_103_b : _GEN_17082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17084 = 9'h68 == r_count_42_io_out ? io_r_104_b : _GEN_17083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17085 = 9'h69 == r_count_42_io_out ? io_r_105_b : _GEN_17084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17086 = 9'h6a == r_count_42_io_out ? io_r_106_b : _GEN_17085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17087 = 9'h6b == r_count_42_io_out ? io_r_107_b : _GEN_17086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17088 = 9'h6c == r_count_42_io_out ? io_r_108_b : _GEN_17087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17089 = 9'h6d == r_count_42_io_out ? io_r_109_b : _GEN_17088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17090 = 9'h6e == r_count_42_io_out ? io_r_110_b : _GEN_17089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17091 = 9'h6f == r_count_42_io_out ? io_r_111_b : _GEN_17090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17092 = 9'h70 == r_count_42_io_out ? io_r_112_b : _GEN_17091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17093 = 9'h71 == r_count_42_io_out ? io_r_113_b : _GEN_17092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17094 = 9'h72 == r_count_42_io_out ? io_r_114_b : _GEN_17093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17095 = 9'h73 == r_count_42_io_out ? io_r_115_b : _GEN_17094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17096 = 9'h74 == r_count_42_io_out ? io_r_116_b : _GEN_17095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17097 = 9'h75 == r_count_42_io_out ? io_r_117_b : _GEN_17096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17098 = 9'h76 == r_count_42_io_out ? io_r_118_b : _GEN_17097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17099 = 9'h77 == r_count_42_io_out ? io_r_119_b : _GEN_17098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17100 = 9'h78 == r_count_42_io_out ? io_r_120_b : _GEN_17099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17101 = 9'h79 == r_count_42_io_out ? io_r_121_b : _GEN_17100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17102 = 9'h7a == r_count_42_io_out ? io_r_122_b : _GEN_17101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17103 = 9'h7b == r_count_42_io_out ? io_r_123_b : _GEN_17102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17104 = 9'h7c == r_count_42_io_out ? io_r_124_b : _GEN_17103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17105 = 9'h7d == r_count_42_io_out ? io_r_125_b : _GEN_17104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17106 = 9'h7e == r_count_42_io_out ? io_r_126_b : _GEN_17105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17107 = 9'h7f == r_count_42_io_out ? io_r_127_b : _GEN_17106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17108 = 9'h80 == r_count_42_io_out ? io_r_128_b : _GEN_17107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17109 = 9'h81 == r_count_42_io_out ? io_r_129_b : _GEN_17108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17110 = 9'h82 == r_count_42_io_out ? io_r_130_b : _GEN_17109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17111 = 9'h83 == r_count_42_io_out ? io_r_131_b : _GEN_17110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17112 = 9'h84 == r_count_42_io_out ? io_r_132_b : _GEN_17111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17113 = 9'h85 == r_count_42_io_out ? io_r_133_b : _GEN_17112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17114 = 9'h86 == r_count_42_io_out ? io_r_134_b : _GEN_17113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17115 = 9'h87 == r_count_42_io_out ? io_r_135_b : _GEN_17114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17116 = 9'h88 == r_count_42_io_out ? io_r_136_b : _GEN_17115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17117 = 9'h89 == r_count_42_io_out ? io_r_137_b : _GEN_17116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17118 = 9'h8a == r_count_42_io_out ? io_r_138_b : _GEN_17117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17119 = 9'h8b == r_count_42_io_out ? io_r_139_b : _GEN_17118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17120 = 9'h8c == r_count_42_io_out ? io_r_140_b : _GEN_17119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17121 = 9'h8d == r_count_42_io_out ? io_r_141_b : _GEN_17120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17122 = 9'h8e == r_count_42_io_out ? io_r_142_b : _GEN_17121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17123 = 9'h8f == r_count_42_io_out ? io_r_143_b : _GEN_17122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17124 = 9'h90 == r_count_42_io_out ? io_r_144_b : _GEN_17123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17125 = 9'h91 == r_count_42_io_out ? io_r_145_b : _GEN_17124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17126 = 9'h92 == r_count_42_io_out ? io_r_146_b : _GEN_17125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17127 = 9'h93 == r_count_42_io_out ? io_r_147_b : _GEN_17126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17128 = 9'h94 == r_count_42_io_out ? io_r_148_b : _GEN_17127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17129 = 9'h95 == r_count_42_io_out ? io_r_149_b : _GEN_17128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17130 = 9'h96 == r_count_42_io_out ? io_r_150_b : _GEN_17129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17131 = 9'h97 == r_count_42_io_out ? io_r_151_b : _GEN_17130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17132 = 9'h98 == r_count_42_io_out ? io_r_152_b : _GEN_17131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17133 = 9'h99 == r_count_42_io_out ? io_r_153_b : _GEN_17132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17134 = 9'h9a == r_count_42_io_out ? io_r_154_b : _GEN_17133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17135 = 9'h9b == r_count_42_io_out ? io_r_155_b : _GEN_17134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17136 = 9'h9c == r_count_42_io_out ? io_r_156_b : _GEN_17135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17137 = 9'h9d == r_count_42_io_out ? io_r_157_b : _GEN_17136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17138 = 9'h9e == r_count_42_io_out ? io_r_158_b : _GEN_17137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17139 = 9'h9f == r_count_42_io_out ? io_r_159_b : _GEN_17138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17140 = 9'ha0 == r_count_42_io_out ? io_r_160_b : _GEN_17139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17141 = 9'ha1 == r_count_42_io_out ? io_r_161_b : _GEN_17140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17142 = 9'ha2 == r_count_42_io_out ? io_r_162_b : _GEN_17141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17143 = 9'ha3 == r_count_42_io_out ? io_r_163_b : _GEN_17142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17144 = 9'ha4 == r_count_42_io_out ? io_r_164_b : _GEN_17143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17145 = 9'ha5 == r_count_42_io_out ? io_r_165_b : _GEN_17144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17146 = 9'ha6 == r_count_42_io_out ? io_r_166_b : _GEN_17145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17147 = 9'ha7 == r_count_42_io_out ? io_r_167_b : _GEN_17146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17148 = 9'ha8 == r_count_42_io_out ? io_r_168_b : _GEN_17147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17149 = 9'ha9 == r_count_42_io_out ? io_r_169_b : _GEN_17148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17150 = 9'haa == r_count_42_io_out ? io_r_170_b : _GEN_17149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17151 = 9'hab == r_count_42_io_out ? io_r_171_b : _GEN_17150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17152 = 9'hac == r_count_42_io_out ? io_r_172_b : _GEN_17151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17153 = 9'had == r_count_42_io_out ? io_r_173_b : _GEN_17152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17154 = 9'hae == r_count_42_io_out ? io_r_174_b : _GEN_17153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17155 = 9'haf == r_count_42_io_out ? io_r_175_b : _GEN_17154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17156 = 9'hb0 == r_count_42_io_out ? io_r_176_b : _GEN_17155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17157 = 9'hb1 == r_count_42_io_out ? io_r_177_b : _GEN_17156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17158 = 9'hb2 == r_count_42_io_out ? io_r_178_b : _GEN_17157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17159 = 9'hb3 == r_count_42_io_out ? io_r_179_b : _GEN_17158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17160 = 9'hb4 == r_count_42_io_out ? io_r_180_b : _GEN_17159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17161 = 9'hb5 == r_count_42_io_out ? io_r_181_b : _GEN_17160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17162 = 9'hb6 == r_count_42_io_out ? io_r_182_b : _GEN_17161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17163 = 9'hb7 == r_count_42_io_out ? io_r_183_b : _GEN_17162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17164 = 9'hb8 == r_count_42_io_out ? io_r_184_b : _GEN_17163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17165 = 9'hb9 == r_count_42_io_out ? io_r_185_b : _GEN_17164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17166 = 9'hba == r_count_42_io_out ? io_r_186_b : _GEN_17165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17167 = 9'hbb == r_count_42_io_out ? io_r_187_b : _GEN_17166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17168 = 9'hbc == r_count_42_io_out ? io_r_188_b : _GEN_17167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17169 = 9'hbd == r_count_42_io_out ? io_r_189_b : _GEN_17168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17170 = 9'hbe == r_count_42_io_out ? io_r_190_b : _GEN_17169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17171 = 9'hbf == r_count_42_io_out ? io_r_191_b : _GEN_17170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17172 = 9'hc0 == r_count_42_io_out ? io_r_192_b : _GEN_17171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17173 = 9'hc1 == r_count_42_io_out ? io_r_193_b : _GEN_17172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17174 = 9'hc2 == r_count_42_io_out ? io_r_194_b : _GEN_17173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17175 = 9'hc3 == r_count_42_io_out ? io_r_195_b : _GEN_17174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17176 = 9'hc4 == r_count_42_io_out ? io_r_196_b : _GEN_17175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17177 = 9'hc5 == r_count_42_io_out ? io_r_197_b : _GEN_17176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17178 = 9'hc6 == r_count_42_io_out ? io_r_198_b : _GEN_17177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17179 = 9'hc7 == r_count_42_io_out ? io_r_199_b : _GEN_17178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17180 = 9'hc8 == r_count_42_io_out ? io_r_200_b : _GEN_17179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17181 = 9'hc9 == r_count_42_io_out ? io_r_201_b : _GEN_17180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17182 = 9'hca == r_count_42_io_out ? io_r_202_b : _GEN_17181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17183 = 9'hcb == r_count_42_io_out ? io_r_203_b : _GEN_17182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17184 = 9'hcc == r_count_42_io_out ? io_r_204_b : _GEN_17183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17185 = 9'hcd == r_count_42_io_out ? io_r_205_b : _GEN_17184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17186 = 9'hce == r_count_42_io_out ? io_r_206_b : _GEN_17185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17187 = 9'hcf == r_count_42_io_out ? io_r_207_b : _GEN_17186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17188 = 9'hd0 == r_count_42_io_out ? io_r_208_b : _GEN_17187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17189 = 9'hd1 == r_count_42_io_out ? io_r_209_b : _GEN_17188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17190 = 9'hd2 == r_count_42_io_out ? io_r_210_b : _GEN_17189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17191 = 9'hd3 == r_count_42_io_out ? io_r_211_b : _GEN_17190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17192 = 9'hd4 == r_count_42_io_out ? io_r_212_b : _GEN_17191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17193 = 9'hd5 == r_count_42_io_out ? io_r_213_b : _GEN_17192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17194 = 9'hd6 == r_count_42_io_out ? io_r_214_b : _GEN_17193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17195 = 9'hd7 == r_count_42_io_out ? io_r_215_b : _GEN_17194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17196 = 9'hd8 == r_count_42_io_out ? io_r_216_b : _GEN_17195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17197 = 9'hd9 == r_count_42_io_out ? io_r_217_b : _GEN_17196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17198 = 9'hda == r_count_42_io_out ? io_r_218_b : _GEN_17197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17199 = 9'hdb == r_count_42_io_out ? io_r_219_b : _GEN_17198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17200 = 9'hdc == r_count_42_io_out ? io_r_220_b : _GEN_17199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17201 = 9'hdd == r_count_42_io_out ? io_r_221_b : _GEN_17200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17202 = 9'hde == r_count_42_io_out ? io_r_222_b : _GEN_17201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17203 = 9'hdf == r_count_42_io_out ? io_r_223_b : _GEN_17202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17204 = 9'he0 == r_count_42_io_out ? io_r_224_b : _GEN_17203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17205 = 9'he1 == r_count_42_io_out ? io_r_225_b : _GEN_17204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17206 = 9'he2 == r_count_42_io_out ? io_r_226_b : _GEN_17205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17207 = 9'he3 == r_count_42_io_out ? io_r_227_b : _GEN_17206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17208 = 9'he4 == r_count_42_io_out ? io_r_228_b : _GEN_17207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17209 = 9'he5 == r_count_42_io_out ? io_r_229_b : _GEN_17208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17210 = 9'he6 == r_count_42_io_out ? io_r_230_b : _GEN_17209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17211 = 9'he7 == r_count_42_io_out ? io_r_231_b : _GEN_17210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17212 = 9'he8 == r_count_42_io_out ? io_r_232_b : _GEN_17211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17213 = 9'he9 == r_count_42_io_out ? io_r_233_b : _GEN_17212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17214 = 9'hea == r_count_42_io_out ? io_r_234_b : _GEN_17213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17215 = 9'heb == r_count_42_io_out ? io_r_235_b : _GEN_17214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17216 = 9'hec == r_count_42_io_out ? io_r_236_b : _GEN_17215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17217 = 9'hed == r_count_42_io_out ? io_r_237_b : _GEN_17216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17218 = 9'hee == r_count_42_io_out ? io_r_238_b : _GEN_17217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17219 = 9'hef == r_count_42_io_out ? io_r_239_b : _GEN_17218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17220 = 9'hf0 == r_count_42_io_out ? io_r_240_b : _GEN_17219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17221 = 9'hf1 == r_count_42_io_out ? io_r_241_b : _GEN_17220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17222 = 9'hf2 == r_count_42_io_out ? io_r_242_b : _GEN_17221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17223 = 9'hf3 == r_count_42_io_out ? io_r_243_b : _GEN_17222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17224 = 9'hf4 == r_count_42_io_out ? io_r_244_b : _GEN_17223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17225 = 9'hf5 == r_count_42_io_out ? io_r_245_b : _GEN_17224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17226 = 9'hf6 == r_count_42_io_out ? io_r_246_b : _GEN_17225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17227 = 9'hf7 == r_count_42_io_out ? io_r_247_b : _GEN_17226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17228 = 9'hf8 == r_count_42_io_out ? io_r_248_b : _GEN_17227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17229 = 9'hf9 == r_count_42_io_out ? io_r_249_b : _GEN_17228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17230 = 9'hfa == r_count_42_io_out ? io_r_250_b : _GEN_17229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17231 = 9'hfb == r_count_42_io_out ? io_r_251_b : _GEN_17230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17232 = 9'hfc == r_count_42_io_out ? io_r_252_b : _GEN_17231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17233 = 9'hfd == r_count_42_io_out ? io_r_253_b : _GEN_17232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17234 = 9'hfe == r_count_42_io_out ? io_r_254_b : _GEN_17233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17235 = 9'hff == r_count_42_io_out ? io_r_255_b : _GEN_17234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17236 = 9'h100 == r_count_42_io_out ? io_r_256_b : _GEN_17235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17237 = 9'h101 == r_count_42_io_out ? io_r_257_b : _GEN_17236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17238 = 9'h102 == r_count_42_io_out ? io_r_258_b : _GEN_17237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17239 = 9'h103 == r_count_42_io_out ? io_r_259_b : _GEN_17238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17240 = 9'h104 == r_count_42_io_out ? io_r_260_b : _GEN_17239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17241 = 9'h105 == r_count_42_io_out ? io_r_261_b : _GEN_17240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17242 = 9'h106 == r_count_42_io_out ? io_r_262_b : _GEN_17241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17243 = 9'h107 == r_count_42_io_out ? io_r_263_b : _GEN_17242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17244 = 9'h108 == r_count_42_io_out ? io_r_264_b : _GEN_17243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17245 = 9'h109 == r_count_42_io_out ? io_r_265_b : _GEN_17244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17246 = 9'h10a == r_count_42_io_out ? io_r_266_b : _GEN_17245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17247 = 9'h10b == r_count_42_io_out ? io_r_267_b : _GEN_17246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17248 = 9'h10c == r_count_42_io_out ? io_r_268_b : _GEN_17247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17249 = 9'h10d == r_count_42_io_out ? io_r_269_b : _GEN_17248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17250 = 9'h10e == r_count_42_io_out ? io_r_270_b : _GEN_17249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17251 = 9'h10f == r_count_42_io_out ? io_r_271_b : _GEN_17250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17252 = 9'h110 == r_count_42_io_out ? io_r_272_b : _GEN_17251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17253 = 9'h111 == r_count_42_io_out ? io_r_273_b : _GEN_17252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17254 = 9'h112 == r_count_42_io_out ? io_r_274_b : _GEN_17253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17255 = 9'h113 == r_count_42_io_out ? io_r_275_b : _GEN_17254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17256 = 9'h114 == r_count_42_io_out ? io_r_276_b : _GEN_17255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17257 = 9'h115 == r_count_42_io_out ? io_r_277_b : _GEN_17256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17258 = 9'h116 == r_count_42_io_out ? io_r_278_b : _GEN_17257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17259 = 9'h117 == r_count_42_io_out ? io_r_279_b : _GEN_17258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17260 = 9'h118 == r_count_42_io_out ? io_r_280_b : _GEN_17259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17261 = 9'h119 == r_count_42_io_out ? io_r_281_b : _GEN_17260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17262 = 9'h11a == r_count_42_io_out ? io_r_282_b : _GEN_17261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17263 = 9'h11b == r_count_42_io_out ? io_r_283_b : _GEN_17262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17264 = 9'h11c == r_count_42_io_out ? io_r_284_b : _GEN_17263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17265 = 9'h11d == r_count_42_io_out ? io_r_285_b : _GEN_17264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17266 = 9'h11e == r_count_42_io_out ? io_r_286_b : _GEN_17265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17267 = 9'h11f == r_count_42_io_out ? io_r_287_b : _GEN_17266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17268 = 9'h120 == r_count_42_io_out ? io_r_288_b : _GEN_17267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17269 = 9'h121 == r_count_42_io_out ? io_r_289_b : _GEN_17268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17270 = 9'h122 == r_count_42_io_out ? io_r_290_b : _GEN_17269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17271 = 9'h123 == r_count_42_io_out ? io_r_291_b : _GEN_17270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17272 = 9'h124 == r_count_42_io_out ? io_r_292_b : _GEN_17271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17273 = 9'h125 == r_count_42_io_out ? io_r_293_b : _GEN_17272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17274 = 9'h126 == r_count_42_io_out ? io_r_294_b : _GEN_17273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17275 = 9'h127 == r_count_42_io_out ? io_r_295_b : _GEN_17274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17276 = 9'h128 == r_count_42_io_out ? io_r_296_b : _GEN_17275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17277 = 9'h129 == r_count_42_io_out ? io_r_297_b : _GEN_17276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17278 = 9'h12a == r_count_42_io_out ? io_r_298_b : _GEN_17277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17279 = 9'h12b == r_count_42_io_out ? io_r_299_b : _GEN_17278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17280 = 9'h12c == r_count_42_io_out ? io_r_300_b : _GEN_17279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17281 = 9'h12d == r_count_42_io_out ? io_r_301_b : _GEN_17280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17282 = 9'h12e == r_count_42_io_out ? io_r_302_b : _GEN_17281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17283 = 9'h12f == r_count_42_io_out ? io_r_303_b : _GEN_17282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17284 = 9'h130 == r_count_42_io_out ? io_r_304_b : _GEN_17283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17285 = 9'h131 == r_count_42_io_out ? io_r_305_b : _GEN_17284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17286 = 9'h132 == r_count_42_io_out ? io_r_306_b : _GEN_17285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17287 = 9'h133 == r_count_42_io_out ? io_r_307_b : _GEN_17286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17288 = 9'h134 == r_count_42_io_out ? io_r_308_b : _GEN_17287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17289 = 9'h135 == r_count_42_io_out ? io_r_309_b : _GEN_17288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17290 = 9'h136 == r_count_42_io_out ? io_r_310_b : _GEN_17289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17291 = 9'h137 == r_count_42_io_out ? io_r_311_b : _GEN_17290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17292 = 9'h138 == r_count_42_io_out ? io_r_312_b : _GEN_17291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17293 = 9'h139 == r_count_42_io_out ? io_r_313_b : _GEN_17292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17294 = 9'h13a == r_count_42_io_out ? io_r_314_b : _GEN_17293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17295 = 9'h13b == r_count_42_io_out ? io_r_315_b : _GEN_17294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17296 = 9'h13c == r_count_42_io_out ? io_r_316_b : _GEN_17295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17297 = 9'h13d == r_count_42_io_out ? io_r_317_b : _GEN_17296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17298 = 9'h13e == r_count_42_io_out ? io_r_318_b : _GEN_17297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17299 = 9'h13f == r_count_42_io_out ? io_r_319_b : _GEN_17298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17300 = 9'h140 == r_count_42_io_out ? io_r_320_b : _GEN_17299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17301 = 9'h141 == r_count_42_io_out ? io_r_321_b : _GEN_17300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17302 = 9'h142 == r_count_42_io_out ? io_r_322_b : _GEN_17301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17303 = 9'h143 == r_count_42_io_out ? io_r_323_b : _GEN_17302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17304 = 9'h144 == r_count_42_io_out ? io_r_324_b : _GEN_17303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17305 = 9'h145 == r_count_42_io_out ? io_r_325_b : _GEN_17304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17306 = 9'h146 == r_count_42_io_out ? io_r_326_b : _GEN_17305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17307 = 9'h147 == r_count_42_io_out ? io_r_327_b : _GEN_17306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17308 = 9'h148 == r_count_42_io_out ? io_r_328_b : _GEN_17307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17309 = 9'h149 == r_count_42_io_out ? io_r_329_b : _GEN_17308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17310 = 9'h14a == r_count_42_io_out ? io_r_330_b : _GEN_17309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17311 = 9'h14b == r_count_42_io_out ? io_r_331_b : _GEN_17310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17312 = 9'h14c == r_count_42_io_out ? io_r_332_b : _GEN_17311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17313 = 9'h14d == r_count_42_io_out ? io_r_333_b : _GEN_17312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17314 = 9'h14e == r_count_42_io_out ? io_r_334_b : _GEN_17313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17315 = 9'h14f == r_count_42_io_out ? io_r_335_b : _GEN_17314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17316 = 9'h150 == r_count_42_io_out ? io_r_336_b : _GEN_17315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17317 = 9'h151 == r_count_42_io_out ? io_r_337_b : _GEN_17316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17318 = 9'h152 == r_count_42_io_out ? io_r_338_b : _GEN_17317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17319 = 9'h153 == r_count_42_io_out ? io_r_339_b : _GEN_17318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17320 = 9'h154 == r_count_42_io_out ? io_r_340_b : _GEN_17319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17321 = 9'h155 == r_count_42_io_out ? io_r_341_b : _GEN_17320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17322 = 9'h156 == r_count_42_io_out ? io_r_342_b : _GEN_17321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17323 = 9'h157 == r_count_42_io_out ? io_r_343_b : _GEN_17322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17324 = 9'h158 == r_count_42_io_out ? io_r_344_b : _GEN_17323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17325 = 9'h159 == r_count_42_io_out ? io_r_345_b : _GEN_17324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17326 = 9'h15a == r_count_42_io_out ? io_r_346_b : _GEN_17325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17327 = 9'h15b == r_count_42_io_out ? io_r_347_b : _GEN_17326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17328 = 9'h15c == r_count_42_io_out ? io_r_348_b : _GEN_17327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17329 = 9'h15d == r_count_42_io_out ? io_r_349_b : _GEN_17328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17330 = 9'h15e == r_count_42_io_out ? io_r_350_b : _GEN_17329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17331 = 9'h15f == r_count_42_io_out ? io_r_351_b : _GEN_17330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17332 = 9'h160 == r_count_42_io_out ? io_r_352_b : _GEN_17331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17333 = 9'h161 == r_count_42_io_out ? io_r_353_b : _GEN_17332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17334 = 9'h162 == r_count_42_io_out ? io_r_354_b : _GEN_17333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17335 = 9'h163 == r_count_42_io_out ? io_r_355_b : _GEN_17334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17336 = 9'h164 == r_count_42_io_out ? io_r_356_b : _GEN_17335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17337 = 9'h165 == r_count_42_io_out ? io_r_357_b : _GEN_17336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17338 = 9'h166 == r_count_42_io_out ? io_r_358_b : _GEN_17337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17339 = 9'h167 == r_count_42_io_out ? io_r_359_b : _GEN_17338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17340 = 9'h168 == r_count_42_io_out ? io_r_360_b : _GEN_17339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17341 = 9'h169 == r_count_42_io_out ? io_r_361_b : _GEN_17340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17342 = 9'h16a == r_count_42_io_out ? io_r_362_b : _GEN_17341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17343 = 9'h16b == r_count_42_io_out ? io_r_363_b : _GEN_17342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17344 = 9'h16c == r_count_42_io_out ? io_r_364_b : _GEN_17343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17345 = 9'h16d == r_count_42_io_out ? io_r_365_b : _GEN_17344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17346 = 9'h16e == r_count_42_io_out ? io_r_366_b : _GEN_17345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17347 = 9'h16f == r_count_42_io_out ? io_r_367_b : _GEN_17346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17348 = 9'h170 == r_count_42_io_out ? io_r_368_b : _GEN_17347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17349 = 9'h171 == r_count_42_io_out ? io_r_369_b : _GEN_17348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17350 = 9'h172 == r_count_42_io_out ? io_r_370_b : _GEN_17349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17351 = 9'h173 == r_count_42_io_out ? io_r_371_b : _GEN_17350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17352 = 9'h174 == r_count_42_io_out ? io_r_372_b : _GEN_17351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17353 = 9'h175 == r_count_42_io_out ? io_r_373_b : _GEN_17352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17354 = 9'h176 == r_count_42_io_out ? io_r_374_b : _GEN_17353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17355 = 9'h177 == r_count_42_io_out ? io_r_375_b : _GEN_17354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17356 = 9'h178 == r_count_42_io_out ? io_r_376_b : _GEN_17355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17357 = 9'h179 == r_count_42_io_out ? io_r_377_b : _GEN_17356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17358 = 9'h17a == r_count_42_io_out ? io_r_378_b : _GEN_17357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17359 = 9'h17b == r_count_42_io_out ? io_r_379_b : _GEN_17358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17360 = 9'h17c == r_count_42_io_out ? io_r_380_b : _GEN_17359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17361 = 9'h17d == r_count_42_io_out ? io_r_381_b : _GEN_17360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17362 = 9'h17e == r_count_42_io_out ? io_r_382_b : _GEN_17361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17363 = 9'h17f == r_count_42_io_out ? io_r_383_b : _GEN_17362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17364 = 9'h180 == r_count_42_io_out ? io_r_384_b : _GEN_17363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17365 = 9'h181 == r_count_42_io_out ? io_r_385_b : _GEN_17364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17366 = 9'h182 == r_count_42_io_out ? io_r_386_b : _GEN_17365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17367 = 9'h183 == r_count_42_io_out ? io_r_387_b : _GEN_17366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17368 = 9'h184 == r_count_42_io_out ? io_r_388_b : _GEN_17367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17369 = 9'h185 == r_count_42_io_out ? io_r_389_b : _GEN_17368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17370 = 9'h186 == r_count_42_io_out ? io_r_390_b : _GEN_17369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17371 = 9'h187 == r_count_42_io_out ? io_r_391_b : _GEN_17370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17372 = 9'h188 == r_count_42_io_out ? io_r_392_b : _GEN_17371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17373 = 9'h189 == r_count_42_io_out ? io_r_393_b : _GEN_17372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17374 = 9'h18a == r_count_42_io_out ? io_r_394_b : _GEN_17373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17375 = 9'h18b == r_count_42_io_out ? io_r_395_b : _GEN_17374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17376 = 9'h18c == r_count_42_io_out ? io_r_396_b : _GEN_17375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17377 = 9'h18d == r_count_42_io_out ? io_r_397_b : _GEN_17376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17378 = 9'h18e == r_count_42_io_out ? io_r_398_b : _GEN_17377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17381 = 9'h1 == r_count_43_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17382 = 9'h2 == r_count_43_io_out ? io_r_2_b : _GEN_17381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17383 = 9'h3 == r_count_43_io_out ? io_r_3_b : _GEN_17382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17384 = 9'h4 == r_count_43_io_out ? io_r_4_b : _GEN_17383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17385 = 9'h5 == r_count_43_io_out ? io_r_5_b : _GEN_17384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17386 = 9'h6 == r_count_43_io_out ? io_r_6_b : _GEN_17385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17387 = 9'h7 == r_count_43_io_out ? io_r_7_b : _GEN_17386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17388 = 9'h8 == r_count_43_io_out ? io_r_8_b : _GEN_17387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17389 = 9'h9 == r_count_43_io_out ? io_r_9_b : _GEN_17388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17390 = 9'ha == r_count_43_io_out ? io_r_10_b : _GEN_17389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17391 = 9'hb == r_count_43_io_out ? io_r_11_b : _GEN_17390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17392 = 9'hc == r_count_43_io_out ? io_r_12_b : _GEN_17391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17393 = 9'hd == r_count_43_io_out ? io_r_13_b : _GEN_17392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17394 = 9'he == r_count_43_io_out ? io_r_14_b : _GEN_17393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17395 = 9'hf == r_count_43_io_out ? io_r_15_b : _GEN_17394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17396 = 9'h10 == r_count_43_io_out ? io_r_16_b : _GEN_17395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17397 = 9'h11 == r_count_43_io_out ? io_r_17_b : _GEN_17396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17398 = 9'h12 == r_count_43_io_out ? io_r_18_b : _GEN_17397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17399 = 9'h13 == r_count_43_io_out ? io_r_19_b : _GEN_17398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17400 = 9'h14 == r_count_43_io_out ? io_r_20_b : _GEN_17399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17401 = 9'h15 == r_count_43_io_out ? io_r_21_b : _GEN_17400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17402 = 9'h16 == r_count_43_io_out ? io_r_22_b : _GEN_17401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17403 = 9'h17 == r_count_43_io_out ? io_r_23_b : _GEN_17402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17404 = 9'h18 == r_count_43_io_out ? io_r_24_b : _GEN_17403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17405 = 9'h19 == r_count_43_io_out ? io_r_25_b : _GEN_17404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17406 = 9'h1a == r_count_43_io_out ? io_r_26_b : _GEN_17405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17407 = 9'h1b == r_count_43_io_out ? io_r_27_b : _GEN_17406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17408 = 9'h1c == r_count_43_io_out ? io_r_28_b : _GEN_17407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17409 = 9'h1d == r_count_43_io_out ? io_r_29_b : _GEN_17408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17410 = 9'h1e == r_count_43_io_out ? io_r_30_b : _GEN_17409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17411 = 9'h1f == r_count_43_io_out ? io_r_31_b : _GEN_17410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17412 = 9'h20 == r_count_43_io_out ? io_r_32_b : _GEN_17411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17413 = 9'h21 == r_count_43_io_out ? io_r_33_b : _GEN_17412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17414 = 9'h22 == r_count_43_io_out ? io_r_34_b : _GEN_17413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17415 = 9'h23 == r_count_43_io_out ? io_r_35_b : _GEN_17414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17416 = 9'h24 == r_count_43_io_out ? io_r_36_b : _GEN_17415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17417 = 9'h25 == r_count_43_io_out ? io_r_37_b : _GEN_17416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17418 = 9'h26 == r_count_43_io_out ? io_r_38_b : _GEN_17417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17419 = 9'h27 == r_count_43_io_out ? io_r_39_b : _GEN_17418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17420 = 9'h28 == r_count_43_io_out ? io_r_40_b : _GEN_17419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17421 = 9'h29 == r_count_43_io_out ? io_r_41_b : _GEN_17420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17422 = 9'h2a == r_count_43_io_out ? io_r_42_b : _GEN_17421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17423 = 9'h2b == r_count_43_io_out ? io_r_43_b : _GEN_17422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17424 = 9'h2c == r_count_43_io_out ? io_r_44_b : _GEN_17423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17425 = 9'h2d == r_count_43_io_out ? io_r_45_b : _GEN_17424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17426 = 9'h2e == r_count_43_io_out ? io_r_46_b : _GEN_17425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17427 = 9'h2f == r_count_43_io_out ? io_r_47_b : _GEN_17426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17428 = 9'h30 == r_count_43_io_out ? io_r_48_b : _GEN_17427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17429 = 9'h31 == r_count_43_io_out ? io_r_49_b : _GEN_17428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17430 = 9'h32 == r_count_43_io_out ? io_r_50_b : _GEN_17429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17431 = 9'h33 == r_count_43_io_out ? io_r_51_b : _GEN_17430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17432 = 9'h34 == r_count_43_io_out ? io_r_52_b : _GEN_17431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17433 = 9'h35 == r_count_43_io_out ? io_r_53_b : _GEN_17432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17434 = 9'h36 == r_count_43_io_out ? io_r_54_b : _GEN_17433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17435 = 9'h37 == r_count_43_io_out ? io_r_55_b : _GEN_17434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17436 = 9'h38 == r_count_43_io_out ? io_r_56_b : _GEN_17435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17437 = 9'h39 == r_count_43_io_out ? io_r_57_b : _GEN_17436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17438 = 9'h3a == r_count_43_io_out ? io_r_58_b : _GEN_17437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17439 = 9'h3b == r_count_43_io_out ? io_r_59_b : _GEN_17438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17440 = 9'h3c == r_count_43_io_out ? io_r_60_b : _GEN_17439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17441 = 9'h3d == r_count_43_io_out ? io_r_61_b : _GEN_17440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17442 = 9'h3e == r_count_43_io_out ? io_r_62_b : _GEN_17441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17443 = 9'h3f == r_count_43_io_out ? io_r_63_b : _GEN_17442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17444 = 9'h40 == r_count_43_io_out ? io_r_64_b : _GEN_17443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17445 = 9'h41 == r_count_43_io_out ? io_r_65_b : _GEN_17444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17446 = 9'h42 == r_count_43_io_out ? io_r_66_b : _GEN_17445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17447 = 9'h43 == r_count_43_io_out ? io_r_67_b : _GEN_17446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17448 = 9'h44 == r_count_43_io_out ? io_r_68_b : _GEN_17447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17449 = 9'h45 == r_count_43_io_out ? io_r_69_b : _GEN_17448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17450 = 9'h46 == r_count_43_io_out ? io_r_70_b : _GEN_17449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17451 = 9'h47 == r_count_43_io_out ? io_r_71_b : _GEN_17450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17452 = 9'h48 == r_count_43_io_out ? io_r_72_b : _GEN_17451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17453 = 9'h49 == r_count_43_io_out ? io_r_73_b : _GEN_17452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17454 = 9'h4a == r_count_43_io_out ? io_r_74_b : _GEN_17453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17455 = 9'h4b == r_count_43_io_out ? io_r_75_b : _GEN_17454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17456 = 9'h4c == r_count_43_io_out ? io_r_76_b : _GEN_17455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17457 = 9'h4d == r_count_43_io_out ? io_r_77_b : _GEN_17456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17458 = 9'h4e == r_count_43_io_out ? io_r_78_b : _GEN_17457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17459 = 9'h4f == r_count_43_io_out ? io_r_79_b : _GEN_17458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17460 = 9'h50 == r_count_43_io_out ? io_r_80_b : _GEN_17459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17461 = 9'h51 == r_count_43_io_out ? io_r_81_b : _GEN_17460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17462 = 9'h52 == r_count_43_io_out ? io_r_82_b : _GEN_17461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17463 = 9'h53 == r_count_43_io_out ? io_r_83_b : _GEN_17462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17464 = 9'h54 == r_count_43_io_out ? io_r_84_b : _GEN_17463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17465 = 9'h55 == r_count_43_io_out ? io_r_85_b : _GEN_17464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17466 = 9'h56 == r_count_43_io_out ? io_r_86_b : _GEN_17465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17467 = 9'h57 == r_count_43_io_out ? io_r_87_b : _GEN_17466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17468 = 9'h58 == r_count_43_io_out ? io_r_88_b : _GEN_17467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17469 = 9'h59 == r_count_43_io_out ? io_r_89_b : _GEN_17468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17470 = 9'h5a == r_count_43_io_out ? io_r_90_b : _GEN_17469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17471 = 9'h5b == r_count_43_io_out ? io_r_91_b : _GEN_17470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17472 = 9'h5c == r_count_43_io_out ? io_r_92_b : _GEN_17471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17473 = 9'h5d == r_count_43_io_out ? io_r_93_b : _GEN_17472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17474 = 9'h5e == r_count_43_io_out ? io_r_94_b : _GEN_17473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17475 = 9'h5f == r_count_43_io_out ? io_r_95_b : _GEN_17474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17476 = 9'h60 == r_count_43_io_out ? io_r_96_b : _GEN_17475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17477 = 9'h61 == r_count_43_io_out ? io_r_97_b : _GEN_17476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17478 = 9'h62 == r_count_43_io_out ? io_r_98_b : _GEN_17477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17479 = 9'h63 == r_count_43_io_out ? io_r_99_b : _GEN_17478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17480 = 9'h64 == r_count_43_io_out ? io_r_100_b : _GEN_17479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17481 = 9'h65 == r_count_43_io_out ? io_r_101_b : _GEN_17480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17482 = 9'h66 == r_count_43_io_out ? io_r_102_b : _GEN_17481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17483 = 9'h67 == r_count_43_io_out ? io_r_103_b : _GEN_17482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17484 = 9'h68 == r_count_43_io_out ? io_r_104_b : _GEN_17483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17485 = 9'h69 == r_count_43_io_out ? io_r_105_b : _GEN_17484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17486 = 9'h6a == r_count_43_io_out ? io_r_106_b : _GEN_17485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17487 = 9'h6b == r_count_43_io_out ? io_r_107_b : _GEN_17486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17488 = 9'h6c == r_count_43_io_out ? io_r_108_b : _GEN_17487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17489 = 9'h6d == r_count_43_io_out ? io_r_109_b : _GEN_17488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17490 = 9'h6e == r_count_43_io_out ? io_r_110_b : _GEN_17489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17491 = 9'h6f == r_count_43_io_out ? io_r_111_b : _GEN_17490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17492 = 9'h70 == r_count_43_io_out ? io_r_112_b : _GEN_17491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17493 = 9'h71 == r_count_43_io_out ? io_r_113_b : _GEN_17492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17494 = 9'h72 == r_count_43_io_out ? io_r_114_b : _GEN_17493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17495 = 9'h73 == r_count_43_io_out ? io_r_115_b : _GEN_17494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17496 = 9'h74 == r_count_43_io_out ? io_r_116_b : _GEN_17495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17497 = 9'h75 == r_count_43_io_out ? io_r_117_b : _GEN_17496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17498 = 9'h76 == r_count_43_io_out ? io_r_118_b : _GEN_17497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17499 = 9'h77 == r_count_43_io_out ? io_r_119_b : _GEN_17498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17500 = 9'h78 == r_count_43_io_out ? io_r_120_b : _GEN_17499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17501 = 9'h79 == r_count_43_io_out ? io_r_121_b : _GEN_17500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17502 = 9'h7a == r_count_43_io_out ? io_r_122_b : _GEN_17501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17503 = 9'h7b == r_count_43_io_out ? io_r_123_b : _GEN_17502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17504 = 9'h7c == r_count_43_io_out ? io_r_124_b : _GEN_17503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17505 = 9'h7d == r_count_43_io_out ? io_r_125_b : _GEN_17504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17506 = 9'h7e == r_count_43_io_out ? io_r_126_b : _GEN_17505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17507 = 9'h7f == r_count_43_io_out ? io_r_127_b : _GEN_17506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17508 = 9'h80 == r_count_43_io_out ? io_r_128_b : _GEN_17507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17509 = 9'h81 == r_count_43_io_out ? io_r_129_b : _GEN_17508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17510 = 9'h82 == r_count_43_io_out ? io_r_130_b : _GEN_17509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17511 = 9'h83 == r_count_43_io_out ? io_r_131_b : _GEN_17510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17512 = 9'h84 == r_count_43_io_out ? io_r_132_b : _GEN_17511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17513 = 9'h85 == r_count_43_io_out ? io_r_133_b : _GEN_17512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17514 = 9'h86 == r_count_43_io_out ? io_r_134_b : _GEN_17513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17515 = 9'h87 == r_count_43_io_out ? io_r_135_b : _GEN_17514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17516 = 9'h88 == r_count_43_io_out ? io_r_136_b : _GEN_17515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17517 = 9'h89 == r_count_43_io_out ? io_r_137_b : _GEN_17516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17518 = 9'h8a == r_count_43_io_out ? io_r_138_b : _GEN_17517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17519 = 9'h8b == r_count_43_io_out ? io_r_139_b : _GEN_17518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17520 = 9'h8c == r_count_43_io_out ? io_r_140_b : _GEN_17519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17521 = 9'h8d == r_count_43_io_out ? io_r_141_b : _GEN_17520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17522 = 9'h8e == r_count_43_io_out ? io_r_142_b : _GEN_17521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17523 = 9'h8f == r_count_43_io_out ? io_r_143_b : _GEN_17522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17524 = 9'h90 == r_count_43_io_out ? io_r_144_b : _GEN_17523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17525 = 9'h91 == r_count_43_io_out ? io_r_145_b : _GEN_17524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17526 = 9'h92 == r_count_43_io_out ? io_r_146_b : _GEN_17525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17527 = 9'h93 == r_count_43_io_out ? io_r_147_b : _GEN_17526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17528 = 9'h94 == r_count_43_io_out ? io_r_148_b : _GEN_17527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17529 = 9'h95 == r_count_43_io_out ? io_r_149_b : _GEN_17528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17530 = 9'h96 == r_count_43_io_out ? io_r_150_b : _GEN_17529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17531 = 9'h97 == r_count_43_io_out ? io_r_151_b : _GEN_17530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17532 = 9'h98 == r_count_43_io_out ? io_r_152_b : _GEN_17531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17533 = 9'h99 == r_count_43_io_out ? io_r_153_b : _GEN_17532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17534 = 9'h9a == r_count_43_io_out ? io_r_154_b : _GEN_17533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17535 = 9'h9b == r_count_43_io_out ? io_r_155_b : _GEN_17534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17536 = 9'h9c == r_count_43_io_out ? io_r_156_b : _GEN_17535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17537 = 9'h9d == r_count_43_io_out ? io_r_157_b : _GEN_17536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17538 = 9'h9e == r_count_43_io_out ? io_r_158_b : _GEN_17537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17539 = 9'h9f == r_count_43_io_out ? io_r_159_b : _GEN_17538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17540 = 9'ha0 == r_count_43_io_out ? io_r_160_b : _GEN_17539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17541 = 9'ha1 == r_count_43_io_out ? io_r_161_b : _GEN_17540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17542 = 9'ha2 == r_count_43_io_out ? io_r_162_b : _GEN_17541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17543 = 9'ha3 == r_count_43_io_out ? io_r_163_b : _GEN_17542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17544 = 9'ha4 == r_count_43_io_out ? io_r_164_b : _GEN_17543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17545 = 9'ha5 == r_count_43_io_out ? io_r_165_b : _GEN_17544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17546 = 9'ha6 == r_count_43_io_out ? io_r_166_b : _GEN_17545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17547 = 9'ha7 == r_count_43_io_out ? io_r_167_b : _GEN_17546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17548 = 9'ha8 == r_count_43_io_out ? io_r_168_b : _GEN_17547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17549 = 9'ha9 == r_count_43_io_out ? io_r_169_b : _GEN_17548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17550 = 9'haa == r_count_43_io_out ? io_r_170_b : _GEN_17549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17551 = 9'hab == r_count_43_io_out ? io_r_171_b : _GEN_17550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17552 = 9'hac == r_count_43_io_out ? io_r_172_b : _GEN_17551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17553 = 9'had == r_count_43_io_out ? io_r_173_b : _GEN_17552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17554 = 9'hae == r_count_43_io_out ? io_r_174_b : _GEN_17553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17555 = 9'haf == r_count_43_io_out ? io_r_175_b : _GEN_17554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17556 = 9'hb0 == r_count_43_io_out ? io_r_176_b : _GEN_17555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17557 = 9'hb1 == r_count_43_io_out ? io_r_177_b : _GEN_17556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17558 = 9'hb2 == r_count_43_io_out ? io_r_178_b : _GEN_17557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17559 = 9'hb3 == r_count_43_io_out ? io_r_179_b : _GEN_17558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17560 = 9'hb4 == r_count_43_io_out ? io_r_180_b : _GEN_17559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17561 = 9'hb5 == r_count_43_io_out ? io_r_181_b : _GEN_17560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17562 = 9'hb6 == r_count_43_io_out ? io_r_182_b : _GEN_17561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17563 = 9'hb7 == r_count_43_io_out ? io_r_183_b : _GEN_17562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17564 = 9'hb8 == r_count_43_io_out ? io_r_184_b : _GEN_17563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17565 = 9'hb9 == r_count_43_io_out ? io_r_185_b : _GEN_17564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17566 = 9'hba == r_count_43_io_out ? io_r_186_b : _GEN_17565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17567 = 9'hbb == r_count_43_io_out ? io_r_187_b : _GEN_17566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17568 = 9'hbc == r_count_43_io_out ? io_r_188_b : _GEN_17567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17569 = 9'hbd == r_count_43_io_out ? io_r_189_b : _GEN_17568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17570 = 9'hbe == r_count_43_io_out ? io_r_190_b : _GEN_17569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17571 = 9'hbf == r_count_43_io_out ? io_r_191_b : _GEN_17570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17572 = 9'hc0 == r_count_43_io_out ? io_r_192_b : _GEN_17571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17573 = 9'hc1 == r_count_43_io_out ? io_r_193_b : _GEN_17572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17574 = 9'hc2 == r_count_43_io_out ? io_r_194_b : _GEN_17573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17575 = 9'hc3 == r_count_43_io_out ? io_r_195_b : _GEN_17574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17576 = 9'hc4 == r_count_43_io_out ? io_r_196_b : _GEN_17575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17577 = 9'hc5 == r_count_43_io_out ? io_r_197_b : _GEN_17576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17578 = 9'hc6 == r_count_43_io_out ? io_r_198_b : _GEN_17577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17579 = 9'hc7 == r_count_43_io_out ? io_r_199_b : _GEN_17578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17580 = 9'hc8 == r_count_43_io_out ? io_r_200_b : _GEN_17579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17581 = 9'hc9 == r_count_43_io_out ? io_r_201_b : _GEN_17580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17582 = 9'hca == r_count_43_io_out ? io_r_202_b : _GEN_17581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17583 = 9'hcb == r_count_43_io_out ? io_r_203_b : _GEN_17582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17584 = 9'hcc == r_count_43_io_out ? io_r_204_b : _GEN_17583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17585 = 9'hcd == r_count_43_io_out ? io_r_205_b : _GEN_17584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17586 = 9'hce == r_count_43_io_out ? io_r_206_b : _GEN_17585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17587 = 9'hcf == r_count_43_io_out ? io_r_207_b : _GEN_17586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17588 = 9'hd0 == r_count_43_io_out ? io_r_208_b : _GEN_17587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17589 = 9'hd1 == r_count_43_io_out ? io_r_209_b : _GEN_17588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17590 = 9'hd2 == r_count_43_io_out ? io_r_210_b : _GEN_17589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17591 = 9'hd3 == r_count_43_io_out ? io_r_211_b : _GEN_17590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17592 = 9'hd4 == r_count_43_io_out ? io_r_212_b : _GEN_17591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17593 = 9'hd5 == r_count_43_io_out ? io_r_213_b : _GEN_17592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17594 = 9'hd6 == r_count_43_io_out ? io_r_214_b : _GEN_17593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17595 = 9'hd7 == r_count_43_io_out ? io_r_215_b : _GEN_17594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17596 = 9'hd8 == r_count_43_io_out ? io_r_216_b : _GEN_17595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17597 = 9'hd9 == r_count_43_io_out ? io_r_217_b : _GEN_17596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17598 = 9'hda == r_count_43_io_out ? io_r_218_b : _GEN_17597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17599 = 9'hdb == r_count_43_io_out ? io_r_219_b : _GEN_17598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17600 = 9'hdc == r_count_43_io_out ? io_r_220_b : _GEN_17599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17601 = 9'hdd == r_count_43_io_out ? io_r_221_b : _GEN_17600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17602 = 9'hde == r_count_43_io_out ? io_r_222_b : _GEN_17601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17603 = 9'hdf == r_count_43_io_out ? io_r_223_b : _GEN_17602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17604 = 9'he0 == r_count_43_io_out ? io_r_224_b : _GEN_17603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17605 = 9'he1 == r_count_43_io_out ? io_r_225_b : _GEN_17604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17606 = 9'he2 == r_count_43_io_out ? io_r_226_b : _GEN_17605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17607 = 9'he3 == r_count_43_io_out ? io_r_227_b : _GEN_17606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17608 = 9'he4 == r_count_43_io_out ? io_r_228_b : _GEN_17607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17609 = 9'he5 == r_count_43_io_out ? io_r_229_b : _GEN_17608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17610 = 9'he6 == r_count_43_io_out ? io_r_230_b : _GEN_17609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17611 = 9'he7 == r_count_43_io_out ? io_r_231_b : _GEN_17610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17612 = 9'he8 == r_count_43_io_out ? io_r_232_b : _GEN_17611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17613 = 9'he9 == r_count_43_io_out ? io_r_233_b : _GEN_17612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17614 = 9'hea == r_count_43_io_out ? io_r_234_b : _GEN_17613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17615 = 9'heb == r_count_43_io_out ? io_r_235_b : _GEN_17614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17616 = 9'hec == r_count_43_io_out ? io_r_236_b : _GEN_17615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17617 = 9'hed == r_count_43_io_out ? io_r_237_b : _GEN_17616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17618 = 9'hee == r_count_43_io_out ? io_r_238_b : _GEN_17617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17619 = 9'hef == r_count_43_io_out ? io_r_239_b : _GEN_17618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17620 = 9'hf0 == r_count_43_io_out ? io_r_240_b : _GEN_17619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17621 = 9'hf1 == r_count_43_io_out ? io_r_241_b : _GEN_17620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17622 = 9'hf2 == r_count_43_io_out ? io_r_242_b : _GEN_17621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17623 = 9'hf3 == r_count_43_io_out ? io_r_243_b : _GEN_17622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17624 = 9'hf4 == r_count_43_io_out ? io_r_244_b : _GEN_17623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17625 = 9'hf5 == r_count_43_io_out ? io_r_245_b : _GEN_17624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17626 = 9'hf6 == r_count_43_io_out ? io_r_246_b : _GEN_17625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17627 = 9'hf7 == r_count_43_io_out ? io_r_247_b : _GEN_17626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17628 = 9'hf8 == r_count_43_io_out ? io_r_248_b : _GEN_17627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17629 = 9'hf9 == r_count_43_io_out ? io_r_249_b : _GEN_17628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17630 = 9'hfa == r_count_43_io_out ? io_r_250_b : _GEN_17629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17631 = 9'hfb == r_count_43_io_out ? io_r_251_b : _GEN_17630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17632 = 9'hfc == r_count_43_io_out ? io_r_252_b : _GEN_17631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17633 = 9'hfd == r_count_43_io_out ? io_r_253_b : _GEN_17632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17634 = 9'hfe == r_count_43_io_out ? io_r_254_b : _GEN_17633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17635 = 9'hff == r_count_43_io_out ? io_r_255_b : _GEN_17634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17636 = 9'h100 == r_count_43_io_out ? io_r_256_b : _GEN_17635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17637 = 9'h101 == r_count_43_io_out ? io_r_257_b : _GEN_17636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17638 = 9'h102 == r_count_43_io_out ? io_r_258_b : _GEN_17637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17639 = 9'h103 == r_count_43_io_out ? io_r_259_b : _GEN_17638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17640 = 9'h104 == r_count_43_io_out ? io_r_260_b : _GEN_17639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17641 = 9'h105 == r_count_43_io_out ? io_r_261_b : _GEN_17640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17642 = 9'h106 == r_count_43_io_out ? io_r_262_b : _GEN_17641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17643 = 9'h107 == r_count_43_io_out ? io_r_263_b : _GEN_17642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17644 = 9'h108 == r_count_43_io_out ? io_r_264_b : _GEN_17643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17645 = 9'h109 == r_count_43_io_out ? io_r_265_b : _GEN_17644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17646 = 9'h10a == r_count_43_io_out ? io_r_266_b : _GEN_17645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17647 = 9'h10b == r_count_43_io_out ? io_r_267_b : _GEN_17646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17648 = 9'h10c == r_count_43_io_out ? io_r_268_b : _GEN_17647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17649 = 9'h10d == r_count_43_io_out ? io_r_269_b : _GEN_17648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17650 = 9'h10e == r_count_43_io_out ? io_r_270_b : _GEN_17649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17651 = 9'h10f == r_count_43_io_out ? io_r_271_b : _GEN_17650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17652 = 9'h110 == r_count_43_io_out ? io_r_272_b : _GEN_17651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17653 = 9'h111 == r_count_43_io_out ? io_r_273_b : _GEN_17652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17654 = 9'h112 == r_count_43_io_out ? io_r_274_b : _GEN_17653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17655 = 9'h113 == r_count_43_io_out ? io_r_275_b : _GEN_17654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17656 = 9'h114 == r_count_43_io_out ? io_r_276_b : _GEN_17655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17657 = 9'h115 == r_count_43_io_out ? io_r_277_b : _GEN_17656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17658 = 9'h116 == r_count_43_io_out ? io_r_278_b : _GEN_17657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17659 = 9'h117 == r_count_43_io_out ? io_r_279_b : _GEN_17658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17660 = 9'h118 == r_count_43_io_out ? io_r_280_b : _GEN_17659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17661 = 9'h119 == r_count_43_io_out ? io_r_281_b : _GEN_17660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17662 = 9'h11a == r_count_43_io_out ? io_r_282_b : _GEN_17661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17663 = 9'h11b == r_count_43_io_out ? io_r_283_b : _GEN_17662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17664 = 9'h11c == r_count_43_io_out ? io_r_284_b : _GEN_17663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17665 = 9'h11d == r_count_43_io_out ? io_r_285_b : _GEN_17664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17666 = 9'h11e == r_count_43_io_out ? io_r_286_b : _GEN_17665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17667 = 9'h11f == r_count_43_io_out ? io_r_287_b : _GEN_17666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17668 = 9'h120 == r_count_43_io_out ? io_r_288_b : _GEN_17667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17669 = 9'h121 == r_count_43_io_out ? io_r_289_b : _GEN_17668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17670 = 9'h122 == r_count_43_io_out ? io_r_290_b : _GEN_17669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17671 = 9'h123 == r_count_43_io_out ? io_r_291_b : _GEN_17670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17672 = 9'h124 == r_count_43_io_out ? io_r_292_b : _GEN_17671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17673 = 9'h125 == r_count_43_io_out ? io_r_293_b : _GEN_17672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17674 = 9'h126 == r_count_43_io_out ? io_r_294_b : _GEN_17673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17675 = 9'h127 == r_count_43_io_out ? io_r_295_b : _GEN_17674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17676 = 9'h128 == r_count_43_io_out ? io_r_296_b : _GEN_17675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17677 = 9'h129 == r_count_43_io_out ? io_r_297_b : _GEN_17676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17678 = 9'h12a == r_count_43_io_out ? io_r_298_b : _GEN_17677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17679 = 9'h12b == r_count_43_io_out ? io_r_299_b : _GEN_17678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17680 = 9'h12c == r_count_43_io_out ? io_r_300_b : _GEN_17679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17681 = 9'h12d == r_count_43_io_out ? io_r_301_b : _GEN_17680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17682 = 9'h12e == r_count_43_io_out ? io_r_302_b : _GEN_17681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17683 = 9'h12f == r_count_43_io_out ? io_r_303_b : _GEN_17682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17684 = 9'h130 == r_count_43_io_out ? io_r_304_b : _GEN_17683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17685 = 9'h131 == r_count_43_io_out ? io_r_305_b : _GEN_17684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17686 = 9'h132 == r_count_43_io_out ? io_r_306_b : _GEN_17685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17687 = 9'h133 == r_count_43_io_out ? io_r_307_b : _GEN_17686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17688 = 9'h134 == r_count_43_io_out ? io_r_308_b : _GEN_17687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17689 = 9'h135 == r_count_43_io_out ? io_r_309_b : _GEN_17688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17690 = 9'h136 == r_count_43_io_out ? io_r_310_b : _GEN_17689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17691 = 9'h137 == r_count_43_io_out ? io_r_311_b : _GEN_17690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17692 = 9'h138 == r_count_43_io_out ? io_r_312_b : _GEN_17691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17693 = 9'h139 == r_count_43_io_out ? io_r_313_b : _GEN_17692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17694 = 9'h13a == r_count_43_io_out ? io_r_314_b : _GEN_17693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17695 = 9'h13b == r_count_43_io_out ? io_r_315_b : _GEN_17694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17696 = 9'h13c == r_count_43_io_out ? io_r_316_b : _GEN_17695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17697 = 9'h13d == r_count_43_io_out ? io_r_317_b : _GEN_17696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17698 = 9'h13e == r_count_43_io_out ? io_r_318_b : _GEN_17697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17699 = 9'h13f == r_count_43_io_out ? io_r_319_b : _GEN_17698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17700 = 9'h140 == r_count_43_io_out ? io_r_320_b : _GEN_17699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17701 = 9'h141 == r_count_43_io_out ? io_r_321_b : _GEN_17700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17702 = 9'h142 == r_count_43_io_out ? io_r_322_b : _GEN_17701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17703 = 9'h143 == r_count_43_io_out ? io_r_323_b : _GEN_17702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17704 = 9'h144 == r_count_43_io_out ? io_r_324_b : _GEN_17703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17705 = 9'h145 == r_count_43_io_out ? io_r_325_b : _GEN_17704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17706 = 9'h146 == r_count_43_io_out ? io_r_326_b : _GEN_17705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17707 = 9'h147 == r_count_43_io_out ? io_r_327_b : _GEN_17706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17708 = 9'h148 == r_count_43_io_out ? io_r_328_b : _GEN_17707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17709 = 9'h149 == r_count_43_io_out ? io_r_329_b : _GEN_17708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17710 = 9'h14a == r_count_43_io_out ? io_r_330_b : _GEN_17709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17711 = 9'h14b == r_count_43_io_out ? io_r_331_b : _GEN_17710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17712 = 9'h14c == r_count_43_io_out ? io_r_332_b : _GEN_17711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17713 = 9'h14d == r_count_43_io_out ? io_r_333_b : _GEN_17712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17714 = 9'h14e == r_count_43_io_out ? io_r_334_b : _GEN_17713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17715 = 9'h14f == r_count_43_io_out ? io_r_335_b : _GEN_17714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17716 = 9'h150 == r_count_43_io_out ? io_r_336_b : _GEN_17715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17717 = 9'h151 == r_count_43_io_out ? io_r_337_b : _GEN_17716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17718 = 9'h152 == r_count_43_io_out ? io_r_338_b : _GEN_17717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17719 = 9'h153 == r_count_43_io_out ? io_r_339_b : _GEN_17718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17720 = 9'h154 == r_count_43_io_out ? io_r_340_b : _GEN_17719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17721 = 9'h155 == r_count_43_io_out ? io_r_341_b : _GEN_17720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17722 = 9'h156 == r_count_43_io_out ? io_r_342_b : _GEN_17721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17723 = 9'h157 == r_count_43_io_out ? io_r_343_b : _GEN_17722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17724 = 9'h158 == r_count_43_io_out ? io_r_344_b : _GEN_17723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17725 = 9'h159 == r_count_43_io_out ? io_r_345_b : _GEN_17724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17726 = 9'h15a == r_count_43_io_out ? io_r_346_b : _GEN_17725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17727 = 9'h15b == r_count_43_io_out ? io_r_347_b : _GEN_17726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17728 = 9'h15c == r_count_43_io_out ? io_r_348_b : _GEN_17727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17729 = 9'h15d == r_count_43_io_out ? io_r_349_b : _GEN_17728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17730 = 9'h15e == r_count_43_io_out ? io_r_350_b : _GEN_17729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17731 = 9'h15f == r_count_43_io_out ? io_r_351_b : _GEN_17730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17732 = 9'h160 == r_count_43_io_out ? io_r_352_b : _GEN_17731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17733 = 9'h161 == r_count_43_io_out ? io_r_353_b : _GEN_17732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17734 = 9'h162 == r_count_43_io_out ? io_r_354_b : _GEN_17733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17735 = 9'h163 == r_count_43_io_out ? io_r_355_b : _GEN_17734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17736 = 9'h164 == r_count_43_io_out ? io_r_356_b : _GEN_17735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17737 = 9'h165 == r_count_43_io_out ? io_r_357_b : _GEN_17736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17738 = 9'h166 == r_count_43_io_out ? io_r_358_b : _GEN_17737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17739 = 9'h167 == r_count_43_io_out ? io_r_359_b : _GEN_17738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17740 = 9'h168 == r_count_43_io_out ? io_r_360_b : _GEN_17739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17741 = 9'h169 == r_count_43_io_out ? io_r_361_b : _GEN_17740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17742 = 9'h16a == r_count_43_io_out ? io_r_362_b : _GEN_17741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17743 = 9'h16b == r_count_43_io_out ? io_r_363_b : _GEN_17742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17744 = 9'h16c == r_count_43_io_out ? io_r_364_b : _GEN_17743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17745 = 9'h16d == r_count_43_io_out ? io_r_365_b : _GEN_17744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17746 = 9'h16e == r_count_43_io_out ? io_r_366_b : _GEN_17745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17747 = 9'h16f == r_count_43_io_out ? io_r_367_b : _GEN_17746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17748 = 9'h170 == r_count_43_io_out ? io_r_368_b : _GEN_17747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17749 = 9'h171 == r_count_43_io_out ? io_r_369_b : _GEN_17748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17750 = 9'h172 == r_count_43_io_out ? io_r_370_b : _GEN_17749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17751 = 9'h173 == r_count_43_io_out ? io_r_371_b : _GEN_17750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17752 = 9'h174 == r_count_43_io_out ? io_r_372_b : _GEN_17751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17753 = 9'h175 == r_count_43_io_out ? io_r_373_b : _GEN_17752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17754 = 9'h176 == r_count_43_io_out ? io_r_374_b : _GEN_17753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17755 = 9'h177 == r_count_43_io_out ? io_r_375_b : _GEN_17754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17756 = 9'h178 == r_count_43_io_out ? io_r_376_b : _GEN_17755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17757 = 9'h179 == r_count_43_io_out ? io_r_377_b : _GEN_17756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17758 = 9'h17a == r_count_43_io_out ? io_r_378_b : _GEN_17757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17759 = 9'h17b == r_count_43_io_out ? io_r_379_b : _GEN_17758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17760 = 9'h17c == r_count_43_io_out ? io_r_380_b : _GEN_17759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17761 = 9'h17d == r_count_43_io_out ? io_r_381_b : _GEN_17760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17762 = 9'h17e == r_count_43_io_out ? io_r_382_b : _GEN_17761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17763 = 9'h17f == r_count_43_io_out ? io_r_383_b : _GEN_17762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17764 = 9'h180 == r_count_43_io_out ? io_r_384_b : _GEN_17763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17765 = 9'h181 == r_count_43_io_out ? io_r_385_b : _GEN_17764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17766 = 9'h182 == r_count_43_io_out ? io_r_386_b : _GEN_17765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17767 = 9'h183 == r_count_43_io_out ? io_r_387_b : _GEN_17766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17768 = 9'h184 == r_count_43_io_out ? io_r_388_b : _GEN_17767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17769 = 9'h185 == r_count_43_io_out ? io_r_389_b : _GEN_17768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17770 = 9'h186 == r_count_43_io_out ? io_r_390_b : _GEN_17769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17771 = 9'h187 == r_count_43_io_out ? io_r_391_b : _GEN_17770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17772 = 9'h188 == r_count_43_io_out ? io_r_392_b : _GEN_17771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17773 = 9'h189 == r_count_43_io_out ? io_r_393_b : _GEN_17772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17774 = 9'h18a == r_count_43_io_out ? io_r_394_b : _GEN_17773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17775 = 9'h18b == r_count_43_io_out ? io_r_395_b : _GEN_17774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17776 = 9'h18c == r_count_43_io_out ? io_r_396_b : _GEN_17775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17777 = 9'h18d == r_count_43_io_out ? io_r_397_b : _GEN_17776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17778 = 9'h18e == r_count_43_io_out ? io_r_398_b : _GEN_17777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17781 = 9'h1 == r_count_44_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17782 = 9'h2 == r_count_44_io_out ? io_r_2_b : _GEN_17781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17783 = 9'h3 == r_count_44_io_out ? io_r_3_b : _GEN_17782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17784 = 9'h4 == r_count_44_io_out ? io_r_4_b : _GEN_17783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17785 = 9'h5 == r_count_44_io_out ? io_r_5_b : _GEN_17784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17786 = 9'h6 == r_count_44_io_out ? io_r_6_b : _GEN_17785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17787 = 9'h7 == r_count_44_io_out ? io_r_7_b : _GEN_17786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17788 = 9'h8 == r_count_44_io_out ? io_r_8_b : _GEN_17787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17789 = 9'h9 == r_count_44_io_out ? io_r_9_b : _GEN_17788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17790 = 9'ha == r_count_44_io_out ? io_r_10_b : _GEN_17789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17791 = 9'hb == r_count_44_io_out ? io_r_11_b : _GEN_17790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17792 = 9'hc == r_count_44_io_out ? io_r_12_b : _GEN_17791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17793 = 9'hd == r_count_44_io_out ? io_r_13_b : _GEN_17792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17794 = 9'he == r_count_44_io_out ? io_r_14_b : _GEN_17793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17795 = 9'hf == r_count_44_io_out ? io_r_15_b : _GEN_17794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17796 = 9'h10 == r_count_44_io_out ? io_r_16_b : _GEN_17795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17797 = 9'h11 == r_count_44_io_out ? io_r_17_b : _GEN_17796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17798 = 9'h12 == r_count_44_io_out ? io_r_18_b : _GEN_17797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17799 = 9'h13 == r_count_44_io_out ? io_r_19_b : _GEN_17798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17800 = 9'h14 == r_count_44_io_out ? io_r_20_b : _GEN_17799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17801 = 9'h15 == r_count_44_io_out ? io_r_21_b : _GEN_17800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17802 = 9'h16 == r_count_44_io_out ? io_r_22_b : _GEN_17801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17803 = 9'h17 == r_count_44_io_out ? io_r_23_b : _GEN_17802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17804 = 9'h18 == r_count_44_io_out ? io_r_24_b : _GEN_17803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17805 = 9'h19 == r_count_44_io_out ? io_r_25_b : _GEN_17804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17806 = 9'h1a == r_count_44_io_out ? io_r_26_b : _GEN_17805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17807 = 9'h1b == r_count_44_io_out ? io_r_27_b : _GEN_17806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17808 = 9'h1c == r_count_44_io_out ? io_r_28_b : _GEN_17807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17809 = 9'h1d == r_count_44_io_out ? io_r_29_b : _GEN_17808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17810 = 9'h1e == r_count_44_io_out ? io_r_30_b : _GEN_17809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17811 = 9'h1f == r_count_44_io_out ? io_r_31_b : _GEN_17810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17812 = 9'h20 == r_count_44_io_out ? io_r_32_b : _GEN_17811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17813 = 9'h21 == r_count_44_io_out ? io_r_33_b : _GEN_17812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17814 = 9'h22 == r_count_44_io_out ? io_r_34_b : _GEN_17813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17815 = 9'h23 == r_count_44_io_out ? io_r_35_b : _GEN_17814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17816 = 9'h24 == r_count_44_io_out ? io_r_36_b : _GEN_17815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17817 = 9'h25 == r_count_44_io_out ? io_r_37_b : _GEN_17816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17818 = 9'h26 == r_count_44_io_out ? io_r_38_b : _GEN_17817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17819 = 9'h27 == r_count_44_io_out ? io_r_39_b : _GEN_17818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17820 = 9'h28 == r_count_44_io_out ? io_r_40_b : _GEN_17819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17821 = 9'h29 == r_count_44_io_out ? io_r_41_b : _GEN_17820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17822 = 9'h2a == r_count_44_io_out ? io_r_42_b : _GEN_17821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17823 = 9'h2b == r_count_44_io_out ? io_r_43_b : _GEN_17822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17824 = 9'h2c == r_count_44_io_out ? io_r_44_b : _GEN_17823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17825 = 9'h2d == r_count_44_io_out ? io_r_45_b : _GEN_17824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17826 = 9'h2e == r_count_44_io_out ? io_r_46_b : _GEN_17825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17827 = 9'h2f == r_count_44_io_out ? io_r_47_b : _GEN_17826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17828 = 9'h30 == r_count_44_io_out ? io_r_48_b : _GEN_17827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17829 = 9'h31 == r_count_44_io_out ? io_r_49_b : _GEN_17828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17830 = 9'h32 == r_count_44_io_out ? io_r_50_b : _GEN_17829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17831 = 9'h33 == r_count_44_io_out ? io_r_51_b : _GEN_17830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17832 = 9'h34 == r_count_44_io_out ? io_r_52_b : _GEN_17831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17833 = 9'h35 == r_count_44_io_out ? io_r_53_b : _GEN_17832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17834 = 9'h36 == r_count_44_io_out ? io_r_54_b : _GEN_17833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17835 = 9'h37 == r_count_44_io_out ? io_r_55_b : _GEN_17834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17836 = 9'h38 == r_count_44_io_out ? io_r_56_b : _GEN_17835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17837 = 9'h39 == r_count_44_io_out ? io_r_57_b : _GEN_17836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17838 = 9'h3a == r_count_44_io_out ? io_r_58_b : _GEN_17837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17839 = 9'h3b == r_count_44_io_out ? io_r_59_b : _GEN_17838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17840 = 9'h3c == r_count_44_io_out ? io_r_60_b : _GEN_17839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17841 = 9'h3d == r_count_44_io_out ? io_r_61_b : _GEN_17840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17842 = 9'h3e == r_count_44_io_out ? io_r_62_b : _GEN_17841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17843 = 9'h3f == r_count_44_io_out ? io_r_63_b : _GEN_17842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17844 = 9'h40 == r_count_44_io_out ? io_r_64_b : _GEN_17843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17845 = 9'h41 == r_count_44_io_out ? io_r_65_b : _GEN_17844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17846 = 9'h42 == r_count_44_io_out ? io_r_66_b : _GEN_17845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17847 = 9'h43 == r_count_44_io_out ? io_r_67_b : _GEN_17846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17848 = 9'h44 == r_count_44_io_out ? io_r_68_b : _GEN_17847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17849 = 9'h45 == r_count_44_io_out ? io_r_69_b : _GEN_17848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17850 = 9'h46 == r_count_44_io_out ? io_r_70_b : _GEN_17849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17851 = 9'h47 == r_count_44_io_out ? io_r_71_b : _GEN_17850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17852 = 9'h48 == r_count_44_io_out ? io_r_72_b : _GEN_17851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17853 = 9'h49 == r_count_44_io_out ? io_r_73_b : _GEN_17852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17854 = 9'h4a == r_count_44_io_out ? io_r_74_b : _GEN_17853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17855 = 9'h4b == r_count_44_io_out ? io_r_75_b : _GEN_17854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17856 = 9'h4c == r_count_44_io_out ? io_r_76_b : _GEN_17855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17857 = 9'h4d == r_count_44_io_out ? io_r_77_b : _GEN_17856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17858 = 9'h4e == r_count_44_io_out ? io_r_78_b : _GEN_17857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17859 = 9'h4f == r_count_44_io_out ? io_r_79_b : _GEN_17858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17860 = 9'h50 == r_count_44_io_out ? io_r_80_b : _GEN_17859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17861 = 9'h51 == r_count_44_io_out ? io_r_81_b : _GEN_17860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17862 = 9'h52 == r_count_44_io_out ? io_r_82_b : _GEN_17861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17863 = 9'h53 == r_count_44_io_out ? io_r_83_b : _GEN_17862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17864 = 9'h54 == r_count_44_io_out ? io_r_84_b : _GEN_17863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17865 = 9'h55 == r_count_44_io_out ? io_r_85_b : _GEN_17864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17866 = 9'h56 == r_count_44_io_out ? io_r_86_b : _GEN_17865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17867 = 9'h57 == r_count_44_io_out ? io_r_87_b : _GEN_17866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17868 = 9'h58 == r_count_44_io_out ? io_r_88_b : _GEN_17867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17869 = 9'h59 == r_count_44_io_out ? io_r_89_b : _GEN_17868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17870 = 9'h5a == r_count_44_io_out ? io_r_90_b : _GEN_17869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17871 = 9'h5b == r_count_44_io_out ? io_r_91_b : _GEN_17870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17872 = 9'h5c == r_count_44_io_out ? io_r_92_b : _GEN_17871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17873 = 9'h5d == r_count_44_io_out ? io_r_93_b : _GEN_17872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17874 = 9'h5e == r_count_44_io_out ? io_r_94_b : _GEN_17873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17875 = 9'h5f == r_count_44_io_out ? io_r_95_b : _GEN_17874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17876 = 9'h60 == r_count_44_io_out ? io_r_96_b : _GEN_17875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17877 = 9'h61 == r_count_44_io_out ? io_r_97_b : _GEN_17876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17878 = 9'h62 == r_count_44_io_out ? io_r_98_b : _GEN_17877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17879 = 9'h63 == r_count_44_io_out ? io_r_99_b : _GEN_17878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17880 = 9'h64 == r_count_44_io_out ? io_r_100_b : _GEN_17879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17881 = 9'h65 == r_count_44_io_out ? io_r_101_b : _GEN_17880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17882 = 9'h66 == r_count_44_io_out ? io_r_102_b : _GEN_17881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17883 = 9'h67 == r_count_44_io_out ? io_r_103_b : _GEN_17882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17884 = 9'h68 == r_count_44_io_out ? io_r_104_b : _GEN_17883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17885 = 9'h69 == r_count_44_io_out ? io_r_105_b : _GEN_17884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17886 = 9'h6a == r_count_44_io_out ? io_r_106_b : _GEN_17885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17887 = 9'h6b == r_count_44_io_out ? io_r_107_b : _GEN_17886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17888 = 9'h6c == r_count_44_io_out ? io_r_108_b : _GEN_17887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17889 = 9'h6d == r_count_44_io_out ? io_r_109_b : _GEN_17888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17890 = 9'h6e == r_count_44_io_out ? io_r_110_b : _GEN_17889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17891 = 9'h6f == r_count_44_io_out ? io_r_111_b : _GEN_17890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17892 = 9'h70 == r_count_44_io_out ? io_r_112_b : _GEN_17891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17893 = 9'h71 == r_count_44_io_out ? io_r_113_b : _GEN_17892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17894 = 9'h72 == r_count_44_io_out ? io_r_114_b : _GEN_17893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17895 = 9'h73 == r_count_44_io_out ? io_r_115_b : _GEN_17894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17896 = 9'h74 == r_count_44_io_out ? io_r_116_b : _GEN_17895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17897 = 9'h75 == r_count_44_io_out ? io_r_117_b : _GEN_17896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17898 = 9'h76 == r_count_44_io_out ? io_r_118_b : _GEN_17897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17899 = 9'h77 == r_count_44_io_out ? io_r_119_b : _GEN_17898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17900 = 9'h78 == r_count_44_io_out ? io_r_120_b : _GEN_17899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17901 = 9'h79 == r_count_44_io_out ? io_r_121_b : _GEN_17900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17902 = 9'h7a == r_count_44_io_out ? io_r_122_b : _GEN_17901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17903 = 9'h7b == r_count_44_io_out ? io_r_123_b : _GEN_17902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17904 = 9'h7c == r_count_44_io_out ? io_r_124_b : _GEN_17903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17905 = 9'h7d == r_count_44_io_out ? io_r_125_b : _GEN_17904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17906 = 9'h7e == r_count_44_io_out ? io_r_126_b : _GEN_17905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17907 = 9'h7f == r_count_44_io_out ? io_r_127_b : _GEN_17906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17908 = 9'h80 == r_count_44_io_out ? io_r_128_b : _GEN_17907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17909 = 9'h81 == r_count_44_io_out ? io_r_129_b : _GEN_17908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17910 = 9'h82 == r_count_44_io_out ? io_r_130_b : _GEN_17909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17911 = 9'h83 == r_count_44_io_out ? io_r_131_b : _GEN_17910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17912 = 9'h84 == r_count_44_io_out ? io_r_132_b : _GEN_17911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17913 = 9'h85 == r_count_44_io_out ? io_r_133_b : _GEN_17912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17914 = 9'h86 == r_count_44_io_out ? io_r_134_b : _GEN_17913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17915 = 9'h87 == r_count_44_io_out ? io_r_135_b : _GEN_17914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17916 = 9'h88 == r_count_44_io_out ? io_r_136_b : _GEN_17915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17917 = 9'h89 == r_count_44_io_out ? io_r_137_b : _GEN_17916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17918 = 9'h8a == r_count_44_io_out ? io_r_138_b : _GEN_17917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17919 = 9'h8b == r_count_44_io_out ? io_r_139_b : _GEN_17918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17920 = 9'h8c == r_count_44_io_out ? io_r_140_b : _GEN_17919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17921 = 9'h8d == r_count_44_io_out ? io_r_141_b : _GEN_17920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17922 = 9'h8e == r_count_44_io_out ? io_r_142_b : _GEN_17921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17923 = 9'h8f == r_count_44_io_out ? io_r_143_b : _GEN_17922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17924 = 9'h90 == r_count_44_io_out ? io_r_144_b : _GEN_17923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17925 = 9'h91 == r_count_44_io_out ? io_r_145_b : _GEN_17924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17926 = 9'h92 == r_count_44_io_out ? io_r_146_b : _GEN_17925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17927 = 9'h93 == r_count_44_io_out ? io_r_147_b : _GEN_17926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17928 = 9'h94 == r_count_44_io_out ? io_r_148_b : _GEN_17927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17929 = 9'h95 == r_count_44_io_out ? io_r_149_b : _GEN_17928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17930 = 9'h96 == r_count_44_io_out ? io_r_150_b : _GEN_17929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17931 = 9'h97 == r_count_44_io_out ? io_r_151_b : _GEN_17930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17932 = 9'h98 == r_count_44_io_out ? io_r_152_b : _GEN_17931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17933 = 9'h99 == r_count_44_io_out ? io_r_153_b : _GEN_17932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17934 = 9'h9a == r_count_44_io_out ? io_r_154_b : _GEN_17933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17935 = 9'h9b == r_count_44_io_out ? io_r_155_b : _GEN_17934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17936 = 9'h9c == r_count_44_io_out ? io_r_156_b : _GEN_17935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17937 = 9'h9d == r_count_44_io_out ? io_r_157_b : _GEN_17936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17938 = 9'h9e == r_count_44_io_out ? io_r_158_b : _GEN_17937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17939 = 9'h9f == r_count_44_io_out ? io_r_159_b : _GEN_17938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17940 = 9'ha0 == r_count_44_io_out ? io_r_160_b : _GEN_17939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17941 = 9'ha1 == r_count_44_io_out ? io_r_161_b : _GEN_17940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17942 = 9'ha2 == r_count_44_io_out ? io_r_162_b : _GEN_17941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17943 = 9'ha3 == r_count_44_io_out ? io_r_163_b : _GEN_17942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17944 = 9'ha4 == r_count_44_io_out ? io_r_164_b : _GEN_17943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17945 = 9'ha5 == r_count_44_io_out ? io_r_165_b : _GEN_17944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17946 = 9'ha6 == r_count_44_io_out ? io_r_166_b : _GEN_17945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17947 = 9'ha7 == r_count_44_io_out ? io_r_167_b : _GEN_17946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17948 = 9'ha8 == r_count_44_io_out ? io_r_168_b : _GEN_17947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17949 = 9'ha9 == r_count_44_io_out ? io_r_169_b : _GEN_17948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17950 = 9'haa == r_count_44_io_out ? io_r_170_b : _GEN_17949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17951 = 9'hab == r_count_44_io_out ? io_r_171_b : _GEN_17950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17952 = 9'hac == r_count_44_io_out ? io_r_172_b : _GEN_17951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17953 = 9'had == r_count_44_io_out ? io_r_173_b : _GEN_17952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17954 = 9'hae == r_count_44_io_out ? io_r_174_b : _GEN_17953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17955 = 9'haf == r_count_44_io_out ? io_r_175_b : _GEN_17954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17956 = 9'hb0 == r_count_44_io_out ? io_r_176_b : _GEN_17955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17957 = 9'hb1 == r_count_44_io_out ? io_r_177_b : _GEN_17956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17958 = 9'hb2 == r_count_44_io_out ? io_r_178_b : _GEN_17957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17959 = 9'hb3 == r_count_44_io_out ? io_r_179_b : _GEN_17958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17960 = 9'hb4 == r_count_44_io_out ? io_r_180_b : _GEN_17959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17961 = 9'hb5 == r_count_44_io_out ? io_r_181_b : _GEN_17960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17962 = 9'hb6 == r_count_44_io_out ? io_r_182_b : _GEN_17961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17963 = 9'hb7 == r_count_44_io_out ? io_r_183_b : _GEN_17962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17964 = 9'hb8 == r_count_44_io_out ? io_r_184_b : _GEN_17963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17965 = 9'hb9 == r_count_44_io_out ? io_r_185_b : _GEN_17964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17966 = 9'hba == r_count_44_io_out ? io_r_186_b : _GEN_17965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17967 = 9'hbb == r_count_44_io_out ? io_r_187_b : _GEN_17966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17968 = 9'hbc == r_count_44_io_out ? io_r_188_b : _GEN_17967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17969 = 9'hbd == r_count_44_io_out ? io_r_189_b : _GEN_17968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17970 = 9'hbe == r_count_44_io_out ? io_r_190_b : _GEN_17969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17971 = 9'hbf == r_count_44_io_out ? io_r_191_b : _GEN_17970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17972 = 9'hc0 == r_count_44_io_out ? io_r_192_b : _GEN_17971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17973 = 9'hc1 == r_count_44_io_out ? io_r_193_b : _GEN_17972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17974 = 9'hc2 == r_count_44_io_out ? io_r_194_b : _GEN_17973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17975 = 9'hc3 == r_count_44_io_out ? io_r_195_b : _GEN_17974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17976 = 9'hc4 == r_count_44_io_out ? io_r_196_b : _GEN_17975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17977 = 9'hc5 == r_count_44_io_out ? io_r_197_b : _GEN_17976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17978 = 9'hc6 == r_count_44_io_out ? io_r_198_b : _GEN_17977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17979 = 9'hc7 == r_count_44_io_out ? io_r_199_b : _GEN_17978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17980 = 9'hc8 == r_count_44_io_out ? io_r_200_b : _GEN_17979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17981 = 9'hc9 == r_count_44_io_out ? io_r_201_b : _GEN_17980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17982 = 9'hca == r_count_44_io_out ? io_r_202_b : _GEN_17981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17983 = 9'hcb == r_count_44_io_out ? io_r_203_b : _GEN_17982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17984 = 9'hcc == r_count_44_io_out ? io_r_204_b : _GEN_17983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17985 = 9'hcd == r_count_44_io_out ? io_r_205_b : _GEN_17984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17986 = 9'hce == r_count_44_io_out ? io_r_206_b : _GEN_17985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17987 = 9'hcf == r_count_44_io_out ? io_r_207_b : _GEN_17986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17988 = 9'hd0 == r_count_44_io_out ? io_r_208_b : _GEN_17987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17989 = 9'hd1 == r_count_44_io_out ? io_r_209_b : _GEN_17988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17990 = 9'hd2 == r_count_44_io_out ? io_r_210_b : _GEN_17989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17991 = 9'hd3 == r_count_44_io_out ? io_r_211_b : _GEN_17990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17992 = 9'hd4 == r_count_44_io_out ? io_r_212_b : _GEN_17991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17993 = 9'hd5 == r_count_44_io_out ? io_r_213_b : _GEN_17992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17994 = 9'hd6 == r_count_44_io_out ? io_r_214_b : _GEN_17993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17995 = 9'hd7 == r_count_44_io_out ? io_r_215_b : _GEN_17994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17996 = 9'hd8 == r_count_44_io_out ? io_r_216_b : _GEN_17995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17997 = 9'hd9 == r_count_44_io_out ? io_r_217_b : _GEN_17996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17998 = 9'hda == r_count_44_io_out ? io_r_218_b : _GEN_17997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17999 = 9'hdb == r_count_44_io_out ? io_r_219_b : _GEN_17998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18000 = 9'hdc == r_count_44_io_out ? io_r_220_b : _GEN_17999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18001 = 9'hdd == r_count_44_io_out ? io_r_221_b : _GEN_18000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18002 = 9'hde == r_count_44_io_out ? io_r_222_b : _GEN_18001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18003 = 9'hdf == r_count_44_io_out ? io_r_223_b : _GEN_18002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18004 = 9'he0 == r_count_44_io_out ? io_r_224_b : _GEN_18003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18005 = 9'he1 == r_count_44_io_out ? io_r_225_b : _GEN_18004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18006 = 9'he2 == r_count_44_io_out ? io_r_226_b : _GEN_18005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18007 = 9'he3 == r_count_44_io_out ? io_r_227_b : _GEN_18006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18008 = 9'he4 == r_count_44_io_out ? io_r_228_b : _GEN_18007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18009 = 9'he5 == r_count_44_io_out ? io_r_229_b : _GEN_18008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18010 = 9'he6 == r_count_44_io_out ? io_r_230_b : _GEN_18009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18011 = 9'he7 == r_count_44_io_out ? io_r_231_b : _GEN_18010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18012 = 9'he8 == r_count_44_io_out ? io_r_232_b : _GEN_18011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18013 = 9'he9 == r_count_44_io_out ? io_r_233_b : _GEN_18012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18014 = 9'hea == r_count_44_io_out ? io_r_234_b : _GEN_18013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18015 = 9'heb == r_count_44_io_out ? io_r_235_b : _GEN_18014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18016 = 9'hec == r_count_44_io_out ? io_r_236_b : _GEN_18015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18017 = 9'hed == r_count_44_io_out ? io_r_237_b : _GEN_18016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18018 = 9'hee == r_count_44_io_out ? io_r_238_b : _GEN_18017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18019 = 9'hef == r_count_44_io_out ? io_r_239_b : _GEN_18018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18020 = 9'hf0 == r_count_44_io_out ? io_r_240_b : _GEN_18019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18021 = 9'hf1 == r_count_44_io_out ? io_r_241_b : _GEN_18020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18022 = 9'hf2 == r_count_44_io_out ? io_r_242_b : _GEN_18021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18023 = 9'hf3 == r_count_44_io_out ? io_r_243_b : _GEN_18022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18024 = 9'hf4 == r_count_44_io_out ? io_r_244_b : _GEN_18023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18025 = 9'hf5 == r_count_44_io_out ? io_r_245_b : _GEN_18024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18026 = 9'hf6 == r_count_44_io_out ? io_r_246_b : _GEN_18025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18027 = 9'hf7 == r_count_44_io_out ? io_r_247_b : _GEN_18026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18028 = 9'hf8 == r_count_44_io_out ? io_r_248_b : _GEN_18027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18029 = 9'hf9 == r_count_44_io_out ? io_r_249_b : _GEN_18028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18030 = 9'hfa == r_count_44_io_out ? io_r_250_b : _GEN_18029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18031 = 9'hfb == r_count_44_io_out ? io_r_251_b : _GEN_18030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18032 = 9'hfc == r_count_44_io_out ? io_r_252_b : _GEN_18031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18033 = 9'hfd == r_count_44_io_out ? io_r_253_b : _GEN_18032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18034 = 9'hfe == r_count_44_io_out ? io_r_254_b : _GEN_18033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18035 = 9'hff == r_count_44_io_out ? io_r_255_b : _GEN_18034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18036 = 9'h100 == r_count_44_io_out ? io_r_256_b : _GEN_18035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18037 = 9'h101 == r_count_44_io_out ? io_r_257_b : _GEN_18036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18038 = 9'h102 == r_count_44_io_out ? io_r_258_b : _GEN_18037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18039 = 9'h103 == r_count_44_io_out ? io_r_259_b : _GEN_18038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18040 = 9'h104 == r_count_44_io_out ? io_r_260_b : _GEN_18039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18041 = 9'h105 == r_count_44_io_out ? io_r_261_b : _GEN_18040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18042 = 9'h106 == r_count_44_io_out ? io_r_262_b : _GEN_18041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18043 = 9'h107 == r_count_44_io_out ? io_r_263_b : _GEN_18042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18044 = 9'h108 == r_count_44_io_out ? io_r_264_b : _GEN_18043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18045 = 9'h109 == r_count_44_io_out ? io_r_265_b : _GEN_18044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18046 = 9'h10a == r_count_44_io_out ? io_r_266_b : _GEN_18045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18047 = 9'h10b == r_count_44_io_out ? io_r_267_b : _GEN_18046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18048 = 9'h10c == r_count_44_io_out ? io_r_268_b : _GEN_18047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18049 = 9'h10d == r_count_44_io_out ? io_r_269_b : _GEN_18048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18050 = 9'h10e == r_count_44_io_out ? io_r_270_b : _GEN_18049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18051 = 9'h10f == r_count_44_io_out ? io_r_271_b : _GEN_18050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18052 = 9'h110 == r_count_44_io_out ? io_r_272_b : _GEN_18051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18053 = 9'h111 == r_count_44_io_out ? io_r_273_b : _GEN_18052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18054 = 9'h112 == r_count_44_io_out ? io_r_274_b : _GEN_18053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18055 = 9'h113 == r_count_44_io_out ? io_r_275_b : _GEN_18054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18056 = 9'h114 == r_count_44_io_out ? io_r_276_b : _GEN_18055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18057 = 9'h115 == r_count_44_io_out ? io_r_277_b : _GEN_18056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18058 = 9'h116 == r_count_44_io_out ? io_r_278_b : _GEN_18057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18059 = 9'h117 == r_count_44_io_out ? io_r_279_b : _GEN_18058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18060 = 9'h118 == r_count_44_io_out ? io_r_280_b : _GEN_18059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18061 = 9'h119 == r_count_44_io_out ? io_r_281_b : _GEN_18060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18062 = 9'h11a == r_count_44_io_out ? io_r_282_b : _GEN_18061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18063 = 9'h11b == r_count_44_io_out ? io_r_283_b : _GEN_18062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18064 = 9'h11c == r_count_44_io_out ? io_r_284_b : _GEN_18063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18065 = 9'h11d == r_count_44_io_out ? io_r_285_b : _GEN_18064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18066 = 9'h11e == r_count_44_io_out ? io_r_286_b : _GEN_18065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18067 = 9'h11f == r_count_44_io_out ? io_r_287_b : _GEN_18066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18068 = 9'h120 == r_count_44_io_out ? io_r_288_b : _GEN_18067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18069 = 9'h121 == r_count_44_io_out ? io_r_289_b : _GEN_18068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18070 = 9'h122 == r_count_44_io_out ? io_r_290_b : _GEN_18069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18071 = 9'h123 == r_count_44_io_out ? io_r_291_b : _GEN_18070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18072 = 9'h124 == r_count_44_io_out ? io_r_292_b : _GEN_18071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18073 = 9'h125 == r_count_44_io_out ? io_r_293_b : _GEN_18072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18074 = 9'h126 == r_count_44_io_out ? io_r_294_b : _GEN_18073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18075 = 9'h127 == r_count_44_io_out ? io_r_295_b : _GEN_18074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18076 = 9'h128 == r_count_44_io_out ? io_r_296_b : _GEN_18075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18077 = 9'h129 == r_count_44_io_out ? io_r_297_b : _GEN_18076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18078 = 9'h12a == r_count_44_io_out ? io_r_298_b : _GEN_18077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18079 = 9'h12b == r_count_44_io_out ? io_r_299_b : _GEN_18078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18080 = 9'h12c == r_count_44_io_out ? io_r_300_b : _GEN_18079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18081 = 9'h12d == r_count_44_io_out ? io_r_301_b : _GEN_18080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18082 = 9'h12e == r_count_44_io_out ? io_r_302_b : _GEN_18081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18083 = 9'h12f == r_count_44_io_out ? io_r_303_b : _GEN_18082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18084 = 9'h130 == r_count_44_io_out ? io_r_304_b : _GEN_18083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18085 = 9'h131 == r_count_44_io_out ? io_r_305_b : _GEN_18084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18086 = 9'h132 == r_count_44_io_out ? io_r_306_b : _GEN_18085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18087 = 9'h133 == r_count_44_io_out ? io_r_307_b : _GEN_18086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18088 = 9'h134 == r_count_44_io_out ? io_r_308_b : _GEN_18087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18089 = 9'h135 == r_count_44_io_out ? io_r_309_b : _GEN_18088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18090 = 9'h136 == r_count_44_io_out ? io_r_310_b : _GEN_18089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18091 = 9'h137 == r_count_44_io_out ? io_r_311_b : _GEN_18090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18092 = 9'h138 == r_count_44_io_out ? io_r_312_b : _GEN_18091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18093 = 9'h139 == r_count_44_io_out ? io_r_313_b : _GEN_18092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18094 = 9'h13a == r_count_44_io_out ? io_r_314_b : _GEN_18093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18095 = 9'h13b == r_count_44_io_out ? io_r_315_b : _GEN_18094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18096 = 9'h13c == r_count_44_io_out ? io_r_316_b : _GEN_18095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18097 = 9'h13d == r_count_44_io_out ? io_r_317_b : _GEN_18096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18098 = 9'h13e == r_count_44_io_out ? io_r_318_b : _GEN_18097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18099 = 9'h13f == r_count_44_io_out ? io_r_319_b : _GEN_18098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18100 = 9'h140 == r_count_44_io_out ? io_r_320_b : _GEN_18099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18101 = 9'h141 == r_count_44_io_out ? io_r_321_b : _GEN_18100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18102 = 9'h142 == r_count_44_io_out ? io_r_322_b : _GEN_18101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18103 = 9'h143 == r_count_44_io_out ? io_r_323_b : _GEN_18102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18104 = 9'h144 == r_count_44_io_out ? io_r_324_b : _GEN_18103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18105 = 9'h145 == r_count_44_io_out ? io_r_325_b : _GEN_18104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18106 = 9'h146 == r_count_44_io_out ? io_r_326_b : _GEN_18105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18107 = 9'h147 == r_count_44_io_out ? io_r_327_b : _GEN_18106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18108 = 9'h148 == r_count_44_io_out ? io_r_328_b : _GEN_18107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18109 = 9'h149 == r_count_44_io_out ? io_r_329_b : _GEN_18108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18110 = 9'h14a == r_count_44_io_out ? io_r_330_b : _GEN_18109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18111 = 9'h14b == r_count_44_io_out ? io_r_331_b : _GEN_18110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18112 = 9'h14c == r_count_44_io_out ? io_r_332_b : _GEN_18111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18113 = 9'h14d == r_count_44_io_out ? io_r_333_b : _GEN_18112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18114 = 9'h14e == r_count_44_io_out ? io_r_334_b : _GEN_18113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18115 = 9'h14f == r_count_44_io_out ? io_r_335_b : _GEN_18114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18116 = 9'h150 == r_count_44_io_out ? io_r_336_b : _GEN_18115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18117 = 9'h151 == r_count_44_io_out ? io_r_337_b : _GEN_18116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18118 = 9'h152 == r_count_44_io_out ? io_r_338_b : _GEN_18117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18119 = 9'h153 == r_count_44_io_out ? io_r_339_b : _GEN_18118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18120 = 9'h154 == r_count_44_io_out ? io_r_340_b : _GEN_18119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18121 = 9'h155 == r_count_44_io_out ? io_r_341_b : _GEN_18120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18122 = 9'h156 == r_count_44_io_out ? io_r_342_b : _GEN_18121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18123 = 9'h157 == r_count_44_io_out ? io_r_343_b : _GEN_18122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18124 = 9'h158 == r_count_44_io_out ? io_r_344_b : _GEN_18123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18125 = 9'h159 == r_count_44_io_out ? io_r_345_b : _GEN_18124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18126 = 9'h15a == r_count_44_io_out ? io_r_346_b : _GEN_18125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18127 = 9'h15b == r_count_44_io_out ? io_r_347_b : _GEN_18126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18128 = 9'h15c == r_count_44_io_out ? io_r_348_b : _GEN_18127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18129 = 9'h15d == r_count_44_io_out ? io_r_349_b : _GEN_18128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18130 = 9'h15e == r_count_44_io_out ? io_r_350_b : _GEN_18129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18131 = 9'h15f == r_count_44_io_out ? io_r_351_b : _GEN_18130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18132 = 9'h160 == r_count_44_io_out ? io_r_352_b : _GEN_18131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18133 = 9'h161 == r_count_44_io_out ? io_r_353_b : _GEN_18132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18134 = 9'h162 == r_count_44_io_out ? io_r_354_b : _GEN_18133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18135 = 9'h163 == r_count_44_io_out ? io_r_355_b : _GEN_18134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18136 = 9'h164 == r_count_44_io_out ? io_r_356_b : _GEN_18135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18137 = 9'h165 == r_count_44_io_out ? io_r_357_b : _GEN_18136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18138 = 9'h166 == r_count_44_io_out ? io_r_358_b : _GEN_18137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18139 = 9'h167 == r_count_44_io_out ? io_r_359_b : _GEN_18138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18140 = 9'h168 == r_count_44_io_out ? io_r_360_b : _GEN_18139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18141 = 9'h169 == r_count_44_io_out ? io_r_361_b : _GEN_18140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18142 = 9'h16a == r_count_44_io_out ? io_r_362_b : _GEN_18141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18143 = 9'h16b == r_count_44_io_out ? io_r_363_b : _GEN_18142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18144 = 9'h16c == r_count_44_io_out ? io_r_364_b : _GEN_18143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18145 = 9'h16d == r_count_44_io_out ? io_r_365_b : _GEN_18144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18146 = 9'h16e == r_count_44_io_out ? io_r_366_b : _GEN_18145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18147 = 9'h16f == r_count_44_io_out ? io_r_367_b : _GEN_18146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18148 = 9'h170 == r_count_44_io_out ? io_r_368_b : _GEN_18147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18149 = 9'h171 == r_count_44_io_out ? io_r_369_b : _GEN_18148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18150 = 9'h172 == r_count_44_io_out ? io_r_370_b : _GEN_18149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18151 = 9'h173 == r_count_44_io_out ? io_r_371_b : _GEN_18150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18152 = 9'h174 == r_count_44_io_out ? io_r_372_b : _GEN_18151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18153 = 9'h175 == r_count_44_io_out ? io_r_373_b : _GEN_18152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18154 = 9'h176 == r_count_44_io_out ? io_r_374_b : _GEN_18153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18155 = 9'h177 == r_count_44_io_out ? io_r_375_b : _GEN_18154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18156 = 9'h178 == r_count_44_io_out ? io_r_376_b : _GEN_18155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18157 = 9'h179 == r_count_44_io_out ? io_r_377_b : _GEN_18156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18158 = 9'h17a == r_count_44_io_out ? io_r_378_b : _GEN_18157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18159 = 9'h17b == r_count_44_io_out ? io_r_379_b : _GEN_18158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18160 = 9'h17c == r_count_44_io_out ? io_r_380_b : _GEN_18159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18161 = 9'h17d == r_count_44_io_out ? io_r_381_b : _GEN_18160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18162 = 9'h17e == r_count_44_io_out ? io_r_382_b : _GEN_18161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18163 = 9'h17f == r_count_44_io_out ? io_r_383_b : _GEN_18162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18164 = 9'h180 == r_count_44_io_out ? io_r_384_b : _GEN_18163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18165 = 9'h181 == r_count_44_io_out ? io_r_385_b : _GEN_18164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18166 = 9'h182 == r_count_44_io_out ? io_r_386_b : _GEN_18165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18167 = 9'h183 == r_count_44_io_out ? io_r_387_b : _GEN_18166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18168 = 9'h184 == r_count_44_io_out ? io_r_388_b : _GEN_18167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18169 = 9'h185 == r_count_44_io_out ? io_r_389_b : _GEN_18168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18170 = 9'h186 == r_count_44_io_out ? io_r_390_b : _GEN_18169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18171 = 9'h187 == r_count_44_io_out ? io_r_391_b : _GEN_18170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18172 = 9'h188 == r_count_44_io_out ? io_r_392_b : _GEN_18171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18173 = 9'h189 == r_count_44_io_out ? io_r_393_b : _GEN_18172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18174 = 9'h18a == r_count_44_io_out ? io_r_394_b : _GEN_18173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18175 = 9'h18b == r_count_44_io_out ? io_r_395_b : _GEN_18174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18176 = 9'h18c == r_count_44_io_out ? io_r_396_b : _GEN_18175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18177 = 9'h18d == r_count_44_io_out ? io_r_397_b : _GEN_18176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18178 = 9'h18e == r_count_44_io_out ? io_r_398_b : _GEN_18177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18181 = 9'h1 == r_count_45_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18182 = 9'h2 == r_count_45_io_out ? io_r_2_b : _GEN_18181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18183 = 9'h3 == r_count_45_io_out ? io_r_3_b : _GEN_18182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18184 = 9'h4 == r_count_45_io_out ? io_r_4_b : _GEN_18183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18185 = 9'h5 == r_count_45_io_out ? io_r_5_b : _GEN_18184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18186 = 9'h6 == r_count_45_io_out ? io_r_6_b : _GEN_18185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18187 = 9'h7 == r_count_45_io_out ? io_r_7_b : _GEN_18186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18188 = 9'h8 == r_count_45_io_out ? io_r_8_b : _GEN_18187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18189 = 9'h9 == r_count_45_io_out ? io_r_9_b : _GEN_18188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18190 = 9'ha == r_count_45_io_out ? io_r_10_b : _GEN_18189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18191 = 9'hb == r_count_45_io_out ? io_r_11_b : _GEN_18190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18192 = 9'hc == r_count_45_io_out ? io_r_12_b : _GEN_18191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18193 = 9'hd == r_count_45_io_out ? io_r_13_b : _GEN_18192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18194 = 9'he == r_count_45_io_out ? io_r_14_b : _GEN_18193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18195 = 9'hf == r_count_45_io_out ? io_r_15_b : _GEN_18194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18196 = 9'h10 == r_count_45_io_out ? io_r_16_b : _GEN_18195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18197 = 9'h11 == r_count_45_io_out ? io_r_17_b : _GEN_18196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18198 = 9'h12 == r_count_45_io_out ? io_r_18_b : _GEN_18197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18199 = 9'h13 == r_count_45_io_out ? io_r_19_b : _GEN_18198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18200 = 9'h14 == r_count_45_io_out ? io_r_20_b : _GEN_18199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18201 = 9'h15 == r_count_45_io_out ? io_r_21_b : _GEN_18200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18202 = 9'h16 == r_count_45_io_out ? io_r_22_b : _GEN_18201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18203 = 9'h17 == r_count_45_io_out ? io_r_23_b : _GEN_18202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18204 = 9'h18 == r_count_45_io_out ? io_r_24_b : _GEN_18203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18205 = 9'h19 == r_count_45_io_out ? io_r_25_b : _GEN_18204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18206 = 9'h1a == r_count_45_io_out ? io_r_26_b : _GEN_18205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18207 = 9'h1b == r_count_45_io_out ? io_r_27_b : _GEN_18206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18208 = 9'h1c == r_count_45_io_out ? io_r_28_b : _GEN_18207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18209 = 9'h1d == r_count_45_io_out ? io_r_29_b : _GEN_18208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18210 = 9'h1e == r_count_45_io_out ? io_r_30_b : _GEN_18209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18211 = 9'h1f == r_count_45_io_out ? io_r_31_b : _GEN_18210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18212 = 9'h20 == r_count_45_io_out ? io_r_32_b : _GEN_18211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18213 = 9'h21 == r_count_45_io_out ? io_r_33_b : _GEN_18212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18214 = 9'h22 == r_count_45_io_out ? io_r_34_b : _GEN_18213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18215 = 9'h23 == r_count_45_io_out ? io_r_35_b : _GEN_18214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18216 = 9'h24 == r_count_45_io_out ? io_r_36_b : _GEN_18215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18217 = 9'h25 == r_count_45_io_out ? io_r_37_b : _GEN_18216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18218 = 9'h26 == r_count_45_io_out ? io_r_38_b : _GEN_18217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18219 = 9'h27 == r_count_45_io_out ? io_r_39_b : _GEN_18218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18220 = 9'h28 == r_count_45_io_out ? io_r_40_b : _GEN_18219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18221 = 9'h29 == r_count_45_io_out ? io_r_41_b : _GEN_18220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18222 = 9'h2a == r_count_45_io_out ? io_r_42_b : _GEN_18221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18223 = 9'h2b == r_count_45_io_out ? io_r_43_b : _GEN_18222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18224 = 9'h2c == r_count_45_io_out ? io_r_44_b : _GEN_18223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18225 = 9'h2d == r_count_45_io_out ? io_r_45_b : _GEN_18224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18226 = 9'h2e == r_count_45_io_out ? io_r_46_b : _GEN_18225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18227 = 9'h2f == r_count_45_io_out ? io_r_47_b : _GEN_18226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18228 = 9'h30 == r_count_45_io_out ? io_r_48_b : _GEN_18227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18229 = 9'h31 == r_count_45_io_out ? io_r_49_b : _GEN_18228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18230 = 9'h32 == r_count_45_io_out ? io_r_50_b : _GEN_18229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18231 = 9'h33 == r_count_45_io_out ? io_r_51_b : _GEN_18230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18232 = 9'h34 == r_count_45_io_out ? io_r_52_b : _GEN_18231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18233 = 9'h35 == r_count_45_io_out ? io_r_53_b : _GEN_18232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18234 = 9'h36 == r_count_45_io_out ? io_r_54_b : _GEN_18233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18235 = 9'h37 == r_count_45_io_out ? io_r_55_b : _GEN_18234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18236 = 9'h38 == r_count_45_io_out ? io_r_56_b : _GEN_18235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18237 = 9'h39 == r_count_45_io_out ? io_r_57_b : _GEN_18236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18238 = 9'h3a == r_count_45_io_out ? io_r_58_b : _GEN_18237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18239 = 9'h3b == r_count_45_io_out ? io_r_59_b : _GEN_18238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18240 = 9'h3c == r_count_45_io_out ? io_r_60_b : _GEN_18239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18241 = 9'h3d == r_count_45_io_out ? io_r_61_b : _GEN_18240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18242 = 9'h3e == r_count_45_io_out ? io_r_62_b : _GEN_18241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18243 = 9'h3f == r_count_45_io_out ? io_r_63_b : _GEN_18242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18244 = 9'h40 == r_count_45_io_out ? io_r_64_b : _GEN_18243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18245 = 9'h41 == r_count_45_io_out ? io_r_65_b : _GEN_18244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18246 = 9'h42 == r_count_45_io_out ? io_r_66_b : _GEN_18245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18247 = 9'h43 == r_count_45_io_out ? io_r_67_b : _GEN_18246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18248 = 9'h44 == r_count_45_io_out ? io_r_68_b : _GEN_18247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18249 = 9'h45 == r_count_45_io_out ? io_r_69_b : _GEN_18248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18250 = 9'h46 == r_count_45_io_out ? io_r_70_b : _GEN_18249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18251 = 9'h47 == r_count_45_io_out ? io_r_71_b : _GEN_18250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18252 = 9'h48 == r_count_45_io_out ? io_r_72_b : _GEN_18251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18253 = 9'h49 == r_count_45_io_out ? io_r_73_b : _GEN_18252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18254 = 9'h4a == r_count_45_io_out ? io_r_74_b : _GEN_18253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18255 = 9'h4b == r_count_45_io_out ? io_r_75_b : _GEN_18254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18256 = 9'h4c == r_count_45_io_out ? io_r_76_b : _GEN_18255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18257 = 9'h4d == r_count_45_io_out ? io_r_77_b : _GEN_18256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18258 = 9'h4e == r_count_45_io_out ? io_r_78_b : _GEN_18257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18259 = 9'h4f == r_count_45_io_out ? io_r_79_b : _GEN_18258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18260 = 9'h50 == r_count_45_io_out ? io_r_80_b : _GEN_18259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18261 = 9'h51 == r_count_45_io_out ? io_r_81_b : _GEN_18260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18262 = 9'h52 == r_count_45_io_out ? io_r_82_b : _GEN_18261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18263 = 9'h53 == r_count_45_io_out ? io_r_83_b : _GEN_18262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18264 = 9'h54 == r_count_45_io_out ? io_r_84_b : _GEN_18263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18265 = 9'h55 == r_count_45_io_out ? io_r_85_b : _GEN_18264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18266 = 9'h56 == r_count_45_io_out ? io_r_86_b : _GEN_18265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18267 = 9'h57 == r_count_45_io_out ? io_r_87_b : _GEN_18266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18268 = 9'h58 == r_count_45_io_out ? io_r_88_b : _GEN_18267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18269 = 9'h59 == r_count_45_io_out ? io_r_89_b : _GEN_18268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18270 = 9'h5a == r_count_45_io_out ? io_r_90_b : _GEN_18269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18271 = 9'h5b == r_count_45_io_out ? io_r_91_b : _GEN_18270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18272 = 9'h5c == r_count_45_io_out ? io_r_92_b : _GEN_18271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18273 = 9'h5d == r_count_45_io_out ? io_r_93_b : _GEN_18272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18274 = 9'h5e == r_count_45_io_out ? io_r_94_b : _GEN_18273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18275 = 9'h5f == r_count_45_io_out ? io_r_95_b : _GEN_18274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18276 = 9'h60 == r_count_45_io_out ? io_r_96_b : _GEN_18275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18277 = 9'h61 == r_count_45_io_out ? io_r_97_b : _GEN_18276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18278 = 9'h62 == r_count_45_io_out ? io_r_98_b : _GEN_18277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18279 = 9'h63 == r_count_45_io_out ? io_r_99_b : _GEN_18278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18280 = 9'h64 == r_count_45_io_out ? io_r_100_b : _GEN_18279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18281 = 9'h65 == r_count_45_io_out ? io_r_101_b : _GEN_18280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18282 = 9'h66 == r_count_45_io_out ? io_r_102_b : _GEN_18281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18283 = 9'h67 == r_count_45_io_out ? io_r_103_b : _GEN_18282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18284 = 9'h68 == r_count_45_io_out ? io_r_104_b : _GEN_18283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18285 = 9'h69 == r_count_45_io_out ? io_r_105_b : _GEN_18284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18286 = 9'h6a == r_count_45_io_out ? io_r_106_b : _GEN_18285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18287 = 9'h6b == r_count_45_io_out ? io_r_107_b : _GEN_18286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18288 = 9'h6c == r_count_45_io_out ? io_r_108_b : _GEN_18287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18289 = 9'h6d == r_count_45_io_out ? io_r_109_b : _GEN_18288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18290 = 9'h6e == r_count_45_io_out ? io_r_110_b : _GEN_18289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18291 = 9'h6f == r_count_45_io_out ? io_r_111_b : _GEN_18290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18292 = 9'h70 == r_count_45_io_out ? io_r_112_b : _GEN_18291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18293 = 9'h71 == r_count_45_io_out ? io_r_113_b : _GEN_18292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18294 = 9'h72 == r_count_45_io_out ? io_r_114_b : _GEN_18293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18295 = 9'h73 == r_count_45_io_out ? io_r_115_b : _GEN_18294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18296 = 9'h74 == r_count_45_io_out ? io_r_116_b : _GEN_18295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18297 = 9'h75 == r_count_45_io_out ? io_r_117_b : _GEN_18296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18298 = 9'h76 == r_count_45_io_out ? io_r_118_b : _GEN_18297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18299 = 9'h77 == r_count_45_io_out ? io_r_119_b : _GEN_18298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18300 = 9'h78 == r_count_45_io_out ? io_r_120_b : _GEN_18299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18301 = 9'h79 == r_count_45_io_out ? io_r_121_b : _GEN_18300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18302 = 9'h7a == r_count_45_io_out ? io_r_122_b : _GEN_18301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18303 = 9'h7b == r_count_45_io_out ? io_r_123_b : _GEN_18302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18304 = 9'h7c == r_count_45_io_out ? io_r_124_b : _GEN_18303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18305 = 9'h7d == r_count_45_io_out ? io_r_125_b : _GEN_18304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18306 = 9'h7e == r_count_45_io_out ? io_r_126_b : _GEN_18305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18307 = 9'h7f == r_count_45_io_out ? io_r_127_b : _GEN_18306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18308 = 9'h80 == r_count_45_io_out ? io_r_128_b : _GEN_18307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18309 = 9'h81 == r_count_45_io_out ? io_r_129_b : _GEN_18308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18310 = 9'h82 == r_count_45_io_out ? io_r_130_b : _GEN_18309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18311 = 9'h83 == r_count_45_io_out ? io_r_131_b : _GEN_18310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18312 = 9'h84 == r_count_45_io_out ? io_r_132_b : _GEN_18311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18313 = 9'h85 == r_count_45_io_out ? io_r_133_b : _GEN_18312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18314 = 9'h86 == r_count_45_io_out ? io_r_134_b : _GEN_18313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18315 = 9'h87 == r_count_45_io_out ? io_r_135_b : _GEN_18314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18316 = 9'h88 == r_count_45_io_out ? io_r_136_b : _GEN_18315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18317 = 9'h89 == r_count_45_io_out ? io_r_137_b : _GEN_18316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18318 = 9'h8a == r_count_45_io_out ? io_r_138_b : _GEN_18317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18319 = 9'h8b == r_count_45_io_out ? io_r_139_b : _GEN_18318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18320 = 9'h8c == r_count_45_io_out ? io_r_140_b : _GEN_18319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18321 = 9'h8d == r_count_45_io_out ? io_r_141_b : _GEN_18320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18322 = 9'h8e == r_count_45_io_out ? io_r_142_b : _GEN_18321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18323 = 9'h8f == r_count_45_io_out ? io_r_143_b : _GEN_18322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18324 = 9'h90 == r_count_45_io_out ? io_r_144_b : _GEN_18323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18325 = 9'h91 == r_count_45_io_out ? io_r_145_b : _GEN_18324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18326 = 9'h92 == r_count_45_io_out ? io_r_146_b : _GEN_18325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18327 = 9'h93 == r_count_45_io_out ? io_r_147_b : _GEN_18326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18328 = 9'h94 == r_count_45_io_out ? io_r_148_b : _GEN_18327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18329 = 9'h95 == r_count_45_io_out ? io_r_149_b : _GEN_18328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18330 = 9'h96 == r_count_45_io_out ? io_r_150_b : _GEN_18329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18331 = 9'h97 == r_count_45_io_out ? io_r_151_b : _GEN_18330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18332 = 9'h98 == r_count_45_io_out ? io_r_152_b : _GEN_18331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18333 = 9'h99 == r_count_45_io_out ? io_r_153_b : _GEN_18332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18334 = 9'h9a == r_count_45_io_out ? io_r_154_b : _GEN_18333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18335 = 9'h9b == r_count_45_io_out ? io_r_155_b : _GEN_18334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18336 = 9'h9c == r_count_45_io_out ? io_r_156_b : _GEN_18335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18337 = 9'h9d == r_count_45_io_out ? io_r_157_b : _GEN_18336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18338 = 9'h9e == r_count_45_io_out ? io_r_158_b : _GEN_18337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18339 = 9'h9f == r_count_45_io_out ? io_r_159_b : _GEN_18338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18340 = 9'ha0 == r_count_45_io_out ? io_r_160_b : _GEN_18339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18341 = 9'ha1 == r_count_45_io_out ? io_r_161_b : _GEN_18340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18342 = 9'ha2 == r_count_45_io_out ? io_r_162_b : _GEN_18341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18343 = 9'ha3 == r_count_45_io_out ? io_r_163_b : _GEN_18342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18344 = 9'ha4 == r_count_45_io_out ? io_r_164_b : _GEN_18343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18345 = 9'ha5 == r_count_45_io_out ? io_r_165_b : _GEN_18344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18346 = 9'ha6 == r_count_45_io_out ? io_r_166_b : _GEN_18345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18347 = 9'ha7 == r_count_45_io_out ? io_r_167_b : _GEN_18346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18348 = 9'ha8 == r_count_45_io_out ? io_r_168_b : _GEN_18347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18349 = 9'ha9 == r_count_45_io_out ? io_r_169_b : _GEN_18348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18350 = 9'haa == r_count_45_io_out ? io_r_170_b : _GEN_18349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18351 = 9'hab == r_count_45_io_out ? io_r_171_b : _GEN_18350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18352 = 9'hac == r_count_45_io_out ? io_r_172_b : _GEN_18351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18353 = 9'had == r_count_45_io_out ? io_r_173_b : _GEN_18352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18354 = 9'hae == r_count_45_io_out ? io_r_174_b : _GEN_18353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18355 = 9'haf == r_count_45_io_out ? io_r_175_b : _GEN_18354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18356 = 9'hb0 == r_count_45_io_out ? io_r_176_b : _GEN_18355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18357 = 9'hb1 == r_count_45_io_out ? io_r_177_b : _GEN_18356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18358 = 9'hb2 == r_count_45_io_out ? io_r_178_b : _GEN_18357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18359 = 9'hb3 == r_count_45_io_out ? io_r_179_b : _GEN_18358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18360 = 9'hb4 == r_count_45_io_out ? io_r_180_b : _GEN_18359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18361 = 9'hb5 == r_count_45_io_out ? io_r_181_b : _GEN_18360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18362 = 9'hb6 == r_count_45_io_out ? io_r_182_b : _GEN_18361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18363 = 9'hb7 == r_count_45_io_out ? io_r_183_b : _GEN_18362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18364 = 9'hb8 == r_count_45_io_out ? io_r_184_b : _GEN_18363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18365 = 9'hb9 == r_count_45_io_out ? io_r_185_b : _GEN_18364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18366 = 9'hba == r_count_45_io_out ? io_r_186_b : _GEN_18365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18367 = 9'hbb == r_count_45_io_out ? io_r_187_b : _GEN_18366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18368 = 9'hbc == r_count_45_io_out ? io_r_188_b : _GEN_18367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18369 = 9'hbd == r_count_45_io_out ? io_r_189_b : _GEN_18368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18370 = 9'hbe == r_count_45_io_out ? io_r_190_b : _GEN_18369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18371 = 9'hbf == r_count_45_io_out ? io_r_191_b : _GEN_18370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18372 = 9'hc0 == r_count_45_io_out ? io_r_192_b : _GEN_18371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18373 = 9'hc1 == r_count_45_io_out ? io_r_193_b : _GEN_18372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18374 = 9'hc2 == r_count_45_io_out ? io_r_194_b : _GEN_18373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18375 = 9'hc3 == r_count_45_io_out ? io_r_195_b : _GEN_18374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18376 = 9'hc4 == r_count_45_io_out ? io_r_196_b : _GEN_18375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18377 = 9'hc5 == r_count_45_io_out ? io_r_197_b : _GEN_18376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18378 = 9'hc6 == r_count_45_io_out ? io_r_198_b : _GEN_18377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18379 = 9'hc7 == r_count_45_io_out ? io_r_199_b : _GEN_18378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18380 = 9'hc8 == r_count_45_io_out ? io_r_200_b : _GEN_18379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18381 = 9'hc9 == r_count_45_io_out ? io_r_201_b : _GEN_18380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18382 = 9'hca == r_count_45_io_out ? io_r_202_b : _GEN_18381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18383 = 9'hcb == r_count_45_io_out ? io_r_203_b : _GEN_18382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18384 = 9'hcc == r_count_45_io_out ? io_r_204_b : _GEN_18383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18385 = 9'hcd == r_count_45_io_out ? io_r_205_b : _GEN_18384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18386 = 9'hce == r_count_45_io_out ? io_r_206_b : _GEN_18385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18387 = 9'hcf == r_count_45_io_out ? io_r_207_b : _GEN_18386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18388 = 9'hd0 == r_count_45_io_out ? io_r_208_b : _GEN_18387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18389 = 9'hd1 == r_count_45_io_out ? io_r_209_b : _GEN_18388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18390 = 9'hd2 == r_count_45_io_out ? io_r_210_b : _GEN_18389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18391 = 9'hd3 == r_count_45_io_out ? io_r_211_b : _GEN_18390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18392 = 9'hd4 == r_count_45_io_out ? io_r_212_b : _GEN_18391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18393 = 9'hd5 == r_count_45_io_out ? io_r_213_b : _GEN_18392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18394 = 9'hd6 == r_count_45_io_out ? io_r_214_b : _GEN_18393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18395 = 9'hd7 == r_count_45_io_out ? io_r_215_b : _GEN_18394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18396 = 9'hd8 == r_count_45_io_out ? io_r_216_b : _GEN_18395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18397 = 9'hd9 == r_count_45_io_out ? io_r_217_b : _GEN_18396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18398 = 9'hda == r_count_45_io_out ? io_r_218_b : _GEN_18397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18399 = 9'hdb == r_count_45_io_out ? io_r_219_b : _GEN_18398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18400 = 9'hdc == r_count_45_io_out ? io_r_220_b : _GEN_18399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18401 = 9'hdd == r_count_45_io_out ? io_r_221_b : _GEN_18400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18402 = 9'hde == r_count_45_io_out ? io_r_222_b : _GEN_18401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18403 = 9'hdf == r_count_45_io_out ? io_r_223_b : _GEN_18402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18404 = 9'he0 == r_count_45_io_out ? io_r_224_b : _GEN_18403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18405 = 9'he1 == r_count_45_io_out ? io_r_225_b : _GEN_18404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18406 = 9'he2 == r_count_45_io_out ? io_r_226_b : _GEN_18405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18407 = 9'he3 == r_count_45_io_out ? io_r_227_b : _GEN_18406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18408 = 9'he4 == r_count_45_io_out ? io_r_228_b : _GEN_18407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18409 = 9'he5 == r_count_45_io_out ? io_r_229_b : _GEN_18408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18410 = 9'he6 == r_count_45_io_out ? io_r_230_b : _GEN_18409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18411 = 9'he7 == r_count_45_io_out ? io_r_231_b : _GEN_18410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18412 = 9'he8 == r_count_45_io_out ? io_r_232_b : _GEN_18411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18413 = 9'he9 == r_count_45_io_out ? io_r_233_b : _GEN_18412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18414 = 9'hea == r_count_45_io_out ? io_r_234_b : _GEN_18413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18415 = 9'heb == r_count_45_io_out ? io_r_235_b : _GEN_18414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18416 = 9'hec == r_count_45_io_out ? io_r_236_b : _GEN_18415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18417 = 9'hed == r_count_45_io_out ? io_r_237_b : _GEN_18416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18418 = 9'hee == r_count_45_io_out ? io_r_238_b : _GEN_18417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18419 = 9'hef == r_count_45_io_out ? io_r_239_b : _GEN_18418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18420 = 9'hf0 == r_count_45_io_out ? io_r_240_b : _GEN_18419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18421 = 9'hf1 == r_count_45_io_out ? io_r_241_b : _GEN_18420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18422 = 9'hf2 == r_count_45_io_out ? io_r_242_b : _GEN_18421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18423 = 9'hf3 == r_count_45_io_out ? io_r_243_b : _GEN_18422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18424 = 9'hf4 == r_count_45_io_out ? io_r_244_b : _GEN_18423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18425 = 9'hf5 == r_count_45_io_out ? io_r_245_b : _GEN_18424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18426 = 9'hf6 == r_count_45_io_out ? io_r_246_b : _GEN_18425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18427 = 9'hf7 == r_count_45_io_out ? io_r_247_b : _GEN_18426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18428 = 9'hf8 == r_count_45_io_out ? io_r_248_b : _GEN_18427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18429 = 9'hf9 == r_count_45_io_out ? io_r_249_b : _GEN_18428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18430 = 9'hfa == r_count_45_io_out ? io_r_250_b : _GEN_18429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18431 = 9'hfb == r_count_45_io_out ? io_r_251_b : _GEN_18430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18432 = 9'hfc == r_count_45_io_out ? io_r_252_b : _GEN_18431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18433 = 9'hfd == r_count_45_io_out ? io_r_253_b : _GEN_18432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18434 = 9'hfe == r_count_45_io_out ? io_r_254_b : _GEN_18433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18435 = 9'hff == r_count_45_io_out ? io_r_255_b : _GEN_18434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18436 = 9'h100 == r_count_45_io_out ? io_r_256_b : _GEN_18435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18437 = 9'h101 == r_count_45_io_out ? io_r_257_b : _GEN_18436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18438 = 9'h102 == r_count_45_io_out ? io_r_258_b : _GEN_18437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18439 = 9'h103 == r_count_45_io_out ? io_r_259_b : _GEN_18438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18440 = 9'h104 == r_count_45_io_out ? io_r_260_b : _GEN_18439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18441 = 9'h105 == r_count_45_io_out ? io_r_261_b : _GEN_18440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18442 = 9'h106 == r_count_45_io_out ? io_r_262_b : _GEN_18441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18443 = 9'h107 == r_count_45_io_out ? io_r_263_b : _GEN_18442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18444 = 9'h108 == r_count_45_io_out ? io_r_264_b : _GEN_18443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18445 = 9'h109 == r_count_45_io_out ? io_r_265_b : _GEN_18444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18446 = 9'h10a == r_count_45_io_out ? io_r_266_b : _GEN_18445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18447 = 9'h10b == r_count_45_io_out ? io_r_267_b : _GEN_18446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18448 = 9'h10c == r_count_45_io_out ? io_r_268_b : _GEN_18447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18449 = 9'h10d == r_count_45_io_out ? io_r_269_b : _GEN_18448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18450 = 9'h10e == r_count_45_io_out ? io_r_270_b : _GEN_18449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18451 = 9'h10f == r_count_45_io_out ? io_r_271_b : _GEN_18450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18452 = 9'h110 == r_count_45_io_out ? io_r_272_b : _GEN_18451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18453 = 9'h111 == r_count_45_io_out ? io_r_273_b : _GEN_18452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18454 = 9'h112 == r_count_45_io_out ? io_r_274_b : _GEN_18453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18455 = 9'h113 == r_count_45_io_out ? io_r_275_b : _GEN_18454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18456 = 9'h114 == r_count_45_io_out ? io_r_276_b : _GEN_18455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18457 = 9'h115 == r_count_45_io_out ? io_r_277_b : _GEN_18456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18458 = 9'h116 == r_count_45_io_out ? io_r_278_b : _GEN_18457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18459 = 9'h117 == r_count_45_io_out ? io_r_279_b : _GEN_18458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18460 = 9'h118 == r_count_45_io_out ? io_r_280_b : _GEN_18459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18461 = 9'h119 == r_count_45_io_out ? io_r_281_b : _GEN_18460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18462 = 9'h11a == r_count_45_io_out ? io_r_282_b : _GEN_18461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18463 = 9'h11b == r_count_45_io_out ? io_r_283_b : _GEN_18462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18464 = 9'h11c == r_count_45_io_out ? io_r_284_b : _GEN_18463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18465 = 9'h11d == r_count_45_io_out ? io_r_285_b : _GEN_18464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18466 = 9'h11e == r_count_45_io_out ? io_r_286_b : _GEN_18465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18467 = 9'h11f == r_count_45_io_out ? io_r_287_b : _GEN_18466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18468 = 9'h120 == r_count_45_io_out ? io_r_288_b : _GEN_18467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18469 = 9'h121 == r_count_45_io_out ? io_r_289_b : _GEN_18468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18470 = 9'h122 == r_count_45_io_out ? io_r_290_b : _GEN_18469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18471 = 9'h123 == r_count_45_io_out ? io_r_291_b : _GEN_18470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18472 = 9'h124 == r_count_45_io_out ? io_r_292_b : _GEN_18471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18473 = 9'h125 == r_count_45_io_out ? io_r_293_b : _GEN_18472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18474 = 9'h126 == r_count_45_io_out ? io_r_294_b : _GEN_18473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18475 = 9'h127 == r_count_45_io_out ? io_r_295_b : _GEN_18474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18476 = 9'h128 == r_count_45_io_out ? io_r_296_b : _GEN_18475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18477 = 9'h129 == r_count_45_io_out ? io_r_297_b : _GEN_18476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18478 = 9'h12a == r_count_45_io_out ? io_r_298_b : _GEN_18477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18479 = 9'h12b == r_count_45_io_out ? io_r_299_b : _GEN_18478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18480 = 9'h12c == r_count_45_io_out ? io_r_300_b : _GEN_18479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18481 = 9'h12d == r_count_45_io_out ? io_r_301_b : _GEN_18480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18482 = 9'h12e == r_count_45_io_out ? io_r_302_b : _GEN_18481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18483 = 9'h12f == r_count_45_io_out ? io_r_303_b : _GEN_18482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18484 = 9'h130 == r_count_45_io_out ? io_r_304_b : _GEN_18483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18485 = 9'h131 == r_count_45_io_out ? io_r_305_b : _GEN_18484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18486 = 9'h132 == r_count_45_io_out ? io_r_306_b : _GEN_18485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18487 = 9'h133 == r_count_45_io_out ? io_r_307_b : _GEN_18486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18488 = 9'h134 == r_count_45_io_out ? io_r_308_b : _GEN_18487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18489 = 9'h135 == r_count_45_io_out ? io_r_309_b : _GEN_18488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18490 = 9'h136 == r_count_45_io_out ? io_r_310_b : _GEN_18489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18491 = 9'h137 == r_count_45_io_out ? io_r_311_b : _GEN_18490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18492 = 9'h138 == r_count_45_io_out ? io_r_312_b : _GEN_18491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18493 = 9'h139 == r_count_45_io_out ? io_r_313_b : _GEN_18492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18494 = 9'h13a == r_count_45_io_out ? io_r_314_b : _GEN_18493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18495 = 9'h13b == r_count_45_io_out ? io_r_315_b : _GEN_18494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18496 = 9'h13c == r_count_45_io_out ? io_r_316_b : _GEN_18495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18497 = 9'h13d == r_count_45_io_out ? io_r_317_b : _GEN_18496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18498 = 9'h13e == r_count_45_io_out ? io_r_318_b : _GEN_18497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18499 = 9'h13f == r_count_45_io_out ? io_r_319_b : _GEN_18498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18500 = 9'h140 == r_count_45_io_out ? io_r_320_b : _GEN_18499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18501 = 9'h141 == r_count_45_io_out ? io_r_321_b : _GEN_18500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18502 = 9'h142 == r_count_45_io_out ? io_r_322_b : _GEN_18501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18503 = 9'h143 == r_count_45_io_out ? io_r_323_b : _GEN_18502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18504 = 9'h144 == r_count_45_io_out ? io_r_324_b : _GEN_18503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18505 = 9'h145 == r_count_45_io_out ? io_r_325_b : _GEN_18504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18506 = 9'h146 == r_count_45_io_out ? io_r_326_b : _GEN_18505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18507 = 9'h147 == r_count_45_io_out ? io_r_327_b : _GEN_18506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18508 = 9'h148 == r_count_45_io_out ? io_r_328_b : _GEN_18507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18509 = 9'h149 == r_count_45_io_out ? io_r_329_b : _GEN_18508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18510 = 9'h14a == r_count_45_io_out ? io_r_330_b : _GEN_18509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18511 = 9'h14b == r_count_45_io_out ? io_r_331_b : _GEN_18510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18512 = 9'h14c == r_count_45_io_out ? io_r_332_b : _GEN_18511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18513 = 9'h14d == r_count_45_io_out ? io_r_333_b : _GEN_18512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18514 = 9'h14e == r_count_45_io_out ? io_r_334_b : _GEN_18513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18515 = 9'h14f == r_count_45_io_out ? io_r_335_b : _GEN_18514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18516 = 9'h150 == r_count_45_io_out ? io_r_336_b : _GEN_18515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18517 = 9'h151 == r_count_45_io_out ? io_r_337_b : _GEN_18516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18518 = 9'h152 == r_count_45_io_out ? io_r_338_b : _GEN_18517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18519 = 9'h153 == r_count_45_io_out ? io_r_339_b : _GEN_18518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18520 = 9'h154 == r_count_45_io_out ? io_r_340_b : _GEN_18519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18521 = 9'h155 == r_count_45_io_out ? io_r_341_b : _GEN_18520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18522 = 9'h156 == r_count_45_io_out ? io_r_342_b : _GEN_18521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18523 = 9'h157 == r_count_45_io_out ? io_r_343_b : _GEN_18522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18524 = 9'h158 == r_count_45_io_out ? io_r_344_b : _GEN_18523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18525 = 9'h159 == r_count_45_io_out ? io_r_345_b : _GEN_18524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18526 = 9'h15a == r_count_45_io_out ? io_r_346_b : _GEN_18525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18527 = 9'h15b == r_count_45_io_out ? io_r_347_b : _GEN_18526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18528 = 9'h15c == r_count_45_io_out ? io_r_348_b : _GEN_18527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18529 = 9'h15d == r_count_45_io_out ? io_r_349_b : _GEN_18528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18530 = 9'h15e == r_count_45_io_out ? io_r_350_b : _GEN_18529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18531 = 9'h15f == r_count_45_io_out ? io_r_351_b : _GEN_18530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18532 = 9'h160 == r_count_45_io_out ? io_r_352_b : _GEN_18531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18533 = 9'h161 == r_count_45_io_out ? io_r_353_b : _GEN_18532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18534 = 9'h162 == r_count_45_io_out ? io_r_354_b : _GEN_18533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18535 = 9'h163 == r_count_45_io_out ? io_r_355_b : _GEN_18534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18536 = 9'h164 == r_count_45_io_out ? io_r_356_b : _GEN_18535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18537 = 9'h165 == r_count_45_io_out ? io_r_357_b : _GEN_18536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18538 = 9'h166 == r_count_45_io_out ? io_r_358_b : _GEN_18537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18539 = 9'h167 == r_count_45_io_out ? io_r_359_b : _GEN_18538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18540 = 9'h168 == r_count_45_io_out ? io_r_360_b : _GEN_18539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18541 = 9'h169 == r_count_45_io_out ? io_r_361_b : _GEN_18540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18542 = 9'h16a == r_count_45_io_out ? io_r_362_b : _GEN_18541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18543 = 9'h16b == r_count_45_io_out ? io_r_363_b : _GEN_18542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18544 = 9'h16c == r_count_45_io_out ? io_r_364_b : _GEN_18543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18545 = 9'h16d == r_count_45_io_out ? io_r_365_b : _GEN_18544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18546 = 9'h16e == r_count_45_io_out ? io_r_366_b : _GEN_18545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18547 = 9'h16f == r_count_45_io_out ? io_r_367_b : _GEN_18546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18548 = 9'h170 == r_count_45_io_out ? io_r_368_b : _GEN_18547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18549 = 9'h171 == r_count_45_io_out ? io_r_369_b : _GEN_18548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18550 = 9'h172 == r_count_45_io_out ? io_r_370_b : _GEN_18549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18551 = 9'h173 == r_count_45_io_out ? io_r_371_b : _GEN_18550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18552 = 9'h174 == r_count_45_io_out ? io_r_372_b : _GEN_18551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18553 = 9'h175 == r_count_45_io_out ? io_r_373_b : _GEN_18552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18554 = 9'h176 == r_count_45_io_out ? io_r_374_b : _GEN_18553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18555 = 9'h177 == r_count_45_io_out ? io_r_375_b : _GEN_18554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18556 = 9'h178 == r_count_45_io_out ? io_r_376_b : _GEN_18555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18557 = 9'h179 == r_count_45_io_out ? io_r_377_b : _GEN_18556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18558 = 9'h17a == r_count_45_io_out ? io_r_378_b : _GEN_18557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18559 = 9'h17b == r_count_45_io_out ? io_r_379_b : _GEN_18558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18560 = 9'h17c == r_count_45_io_out ? io_r_380_b : _GEN_18559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18561 = 9'h17d == r_count_45_io_out ? io_r_381_b : _GEN_18560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18562 = 9'h17e == r_count_45_io_out ? io_r_382_b : _GEN_18561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18563 = 9'h17f == r_count_45_io_out ? io_r_383_b : _GEN_18562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18564 = 9'h180 == r_count_45_io_out ? io_r_384_b : _GEN_18563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18565 = 9'h181 == r_count_45_io_out ? io_r_385_b : _GEN_18564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18566 = 9'h182 == r_count_45_io_out ? io_r_386_b : _GEN_18565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18567 = 9'h183 == r_count_45_io_out ? io_r_387_b : _GEN_18566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18568 = 9'h184 == r_count_45_io_out ? io_r_388_b : _GEN_18567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18569 = 9'h185 == r_count_45_io_out ? io_r_389_b : _GEN_18568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18570 = 9'h186 == r_count_45_io_out ? io_r_390_b : _GEN_18569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18571 = 9'h187 == r_count_45_io_out ? io_r_391_b : _GEN_18570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18572 = 9'h188 == r_count_45_io_out ? io_r_392_b : _GEN_18571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18573 = 9'h189 == r_count_45_io_out ? io_r_393_b : _GEN_18572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18574 = 9'h18a == r_count_45_io_out ? io_r_394_b : _GEN_18573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18575 = 9'h18b == r_count_45_io_out ? io_r_395_b : _GEN_18574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18576 = 9'h18c == r_count_45_io_out ? io_r_396_b : _GEN_18575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18577 = 9'h18d == r_count_45_io_out ? io_r_397_b : _GEN_18576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18578 = 9'h18e == r_count_45_io_out ? io_r_398_b : _GEN_18577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18581 = 9'h1 == r_count_46_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18582 = 9'h2 == r_count_46_io_out ? io_r_2_b : _GEN_18581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18583 = 9'h3 == r_count_46_io_out ? io_r_3_b : _GEN_18582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18584 = 9'h4 == r_count_46_io_out ? io_r_4_b : _GEN_18583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18585 = 9'h5 == r_count_46_io_out ? io_r_5_b : _GEN_18584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18586 = 9'h6 == r_count_46_io_out ? io_r_6_b : _GEN_18585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18587 = 9'h7 == r_count_46_io_out ? io_r_7_b : _GEN_18586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18588 = 9'h8 == r_count_46_io_out ? io_r_8_b : _GEN_18587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18589 = 9'h9 == r_count_46_io_out ? io_r_9_b : _GEN_18588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18590 = 9'ha == r_count_46_io_out ? io_r_10_b : _GEN_18589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18591 = 9'hb == r_count_46_io_out ? io_r_11_b : _GEN_18590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18592 = 9'hc == r_count_46_io_out ? io_r_12_b : _GEN_18591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18593 = 9'hd == r_count_46_io_out ? io_r_13_b : _GEN_18592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18594 = 9'he == r_count_46_io_out ? io_r_14_b : _GEN_18593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18595 = 9'hf == r_count_46_io_out ? io_r_15_b : _GEN_18594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18596 = 9'h10 == r_count_46_io_out ? io_r_16_b : _GEN_18595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18597 = 9'h11 == r_count_46_io_out ? io_r_17_b : _GEN_18596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18598 = 9'h12 == r_count_46_io_out ? io_r_18_b : _GEN_18597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18599 = 9'h13 == r_count_46_io_out ? io_r_19_b : _GEN_18598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18600 = 9'h14 == r_count_46_io_out ? io_r_20_b : _GEN_18599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18601 = 9'h15 == r_count_46_io_out ? io_r_21_b : _GEN_18600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18602 = 9'h16 == r_count_46_io_out ? io_r_22_b : _GEN_18601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18603 = 9'h17 == r_count_46_io_out ? io_r_23_b : _GEN_18602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18604 = 9'h18 == r_count_46_io_out ? io_r_24_b : _GEN_18603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18605 = 9'h19 == r_count_46_io_out ? io_r_25_b : _GEN_18604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18606 = 9'h1a == r_count_46_io_out ? io_r_26_b : _GEN_18605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18607 = 9'h1b == r_count_46_io_out ? io_r_27_b : _GEN_18606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18608 = 9'h1c == r_count_46_io_out ? io_r_28_b : _GEN_18607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18609 = 9'h1d == r_count_46_io_out ? io_r_29_b : _GEN_18608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18610 = 9'h1e == r_count_46_io_out ? io_r_30_b : _GEN_18609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18611 = 9'h1f == r_count_46_io_out ? io_r_31_b : _GEN_18610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18612 = 9'h20 == r_count_46_io_out ? io_r_32_b : _GEN_18611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18613 = 9'h21 == r_count_46_io_out ? io_r_33_b : _GEN_18612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18614 = 9'h22 == r_count_46_io_out ? io_r_34_b : _GEN_18613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18615 = 9'h23 == r_count_46_io_out ? io_r_35_b : _GEN_18614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18616 = 9'h24 == r_count_46_io_out ? io_r_36_b : _GEN_18615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18617 = 9'h25 == r_count_46_io_out ? io_r_37_b : _GEN_18616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18618 = 9'h26 == r_count_46_io_out ? io_r_38_b : _GEN_18617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18619 = 9'h27 == r_count_46_io_out ? io_r_39_b : _GEN_18618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18620 = 9'h28 == r_count_46_io_out ? io_r_40_b : _GEN_18619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18621 = 9'h29 == r_count_46_io_out ? io_r_41_b : _GEN_18620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18622 = 9'h2a == r_count_46_io_out ? io_r_42_b : _GEN_18621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18623 = 9'h2b == r_count_46_io_out ? io_r_43_b : _GEN_18622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18624 = 9'h2c == r_count_46_io_out ? io_r_44_b : _GEN_18623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18625 = 9'h2d == r_count_46_io_out ? io_r_45_b : _GEN_18624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18626 = 9'h2e == r_count_46_io_out ? io_r_46_b : _GEN_18625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18627 = 9'h2f == r_count_46_io_out ? io_r_47_b : _GEN_18626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18628 = 9'h30 == r_count_46_io_out ? io_r_48_b : _GEN_18627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18629 = 9'h31 == r_count_46_io_out ? io_r_49_b : _GEN_18628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18630 = 9'h32 == r_count_46_io_out ? io_r_50_b : _GEN_18629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18631 = 9'h33 == r_count_46_io_out ? io_r_51_b : _GEN_18630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18632 = 9'h34 == r_count_46_io_out ? io_r_52_b : _GEN_18631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18633 = 9'h35 == r_count_46_io_out ? io_r_53_b : _GEN_18632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18634 = 9'h36 == r_count_46_io_out ? io_r_54_b : _GEN_18633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18635 = 9'h37 == r_count_46_io_out ? io_r_55_b : _GEN_18634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18636 = 9'h38 == r_count_46_io_out ? io_r_56_b : _GEN_18635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18637 = 9'h39 == r_count_46_io_out ? io_r_57_b : _GEN_18636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18638 = 9'h3a == r_count_46_io_out ? io_r_58_b : _GEN_18637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18639 = 9'h3b == r_count_46_io_out ? io_r_59_b : _GEN_18638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18640 = 9'h3c == r_count_46_io_out ? io_r_60_b : _GEN_18639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18641 = 9'h3d == r_count_46_io_out ? io_r_61_b : _GEN_18640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18642 = 9'h3e == r_count_46_io_out ? io_r_62_b : _GEN_18641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18643 = 9'h3f == r_count_46_io_out ? io_r_63_b : _GEN_18642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18644 = 9'h40 == r_count_46_io_out ? io_r_64_b : _GEN_18643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18645 = 9'h41 == r_count_46_io_out ? io_r_65_b : _GEN_18644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18646 = 9'h42 == r_count_46_io_out ? io_r_66_b : _GEN_18645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18647 = 9'h43 == r_count_46_io_out ? io_r_67_b : _GEN_18646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18648 = 9'h44 == r_count_46_io_out ? io_r_68_b : _GEN_18647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18649 = 9'h45 == r_count_46_io_out ? io_r_69_b : _GEN_18648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18650 = 9'h46 == r_count_46_io_out ? io_r_70_b : _GEN_18649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18651 = 9'h47 == r_count_46_io_out ? io_r_71_b : _GEN_18650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18652 = 9'h48 == r_count_46_io_out ? io_r_72_b : _GEN_18651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18653 = 9'h49 == r_count_46_io_out ? io_r_73_b : _GEN_18652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18654 = 9'h4a == r_count_46_io_out ? io_r_74_b : _GEN_18653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18655 = 9'h4b == r_count_46_io_out ? io_r_75_b : _GEN_18654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18656 = 9'h4c == r_count_46_io_out ? io_r_76_b : _GEN_18655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18657 = 9'h4d == r_count_46_io_out ? io_r_77_b : _GEN_18656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18658 = 9'h4e == r_count_46_io_out ? io_r_78_b : _GEN_18657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18659 = 9'h4f == r_count_46_io_out ? io_r_79_b : _GEN_18658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18660 = 9'h50 == r_count_46_io_out ? io_r_80_b : _GEN_18659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18661 = 9'h51 == r_count_46_io_out ? io_r_81_b : _GEN_18660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18662 = 9'h52 == r_count_46_io_out ? io_r_82_b : _GEN_18661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18663 = 9'h53 == r_count_46_io_out ? io_r_83_b : _GEN_18662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18664 = 9'h54 == r_count_46_io_out ? io_r_84_b : _GEN_18663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18665 = 9'h55 == r_count_46_io_out ? io_r_85_b : _GEN_18664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18666 = 9'h56 == r_count_46_io_out ? io_r_86_b : _GEN_18665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18667 = 9'h57 == r_count_46_io_out ? io_r_87_b : _GEN_18666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18668 = 9'h58 == r_count_46_io_out ? io_r_88_b : _GEN_18667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18669 = 9'h59 == r_count_46_io_out ? io_r_89_b : _GEN_18668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18670 = 9'h5a == r_count_46_io_out ? io_r_90_b : _GEN_18669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18671 = 9'h5b == r_count_46_io_out ? io_r_91_b : _GEN_18670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18672 = 9'h5c == r_count_46_io_out ? io_r_92_b : _GEN_18671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18673 = 9'h5d == r_count_46_io_out ? io_r_93_b : _GEN_18672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18674 = 9'h5e == r_count_46_io_out ? io_r_94_b : _GEN_18673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18675 = 9'h5f == r_count_46_io_out ? io_r_95_b : _GEN_18674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18676 = 9'h60 == r_count_46_io_out ? io_r_96_b : _GEN_18675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18677 = 9'h61 == r_count_46_io_out ? io_r_97_b : _GEN_18676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18678 = 9'h62 == r_count_46_io_out ? io_r_98_b : _GEN_18677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18679 = 9'h63 == r_count_46_io_out ? io_r_99_b : _GEN_18678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18680 = 9'h64 == r_count_46_io_out ? io_r_100_b : _GEN_18679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18681 = 9'h65 == r_count_46_io_out ? io_r_101_b : _GEN_18680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18682 = 9'h66 == r_count_46_io_out ? io_r_102_b : _GEN_18681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18683 = 9'h67 == r_count_46_io_out ? io_r_103_b : _GEN_18682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18684 = 9'h68 == r_count_46_io_out ? io_r_104_b : _GEN_18683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18685 = 9'h69 == r_count_46_io_out ? io_r_105_b : _GEN_18684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18686 = 9'h6a == r_count_46_io_out ? io_r_106_b : _GEN_18685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18687 = 9'h6b == r_count_46_io_out ? io_r_107_b : _GEN_18686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18688 = 9'h6c == r_count_46_io_out ? io_r_108_b : _GEN_18687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18689 = 9'h6d == r_count_46_io_out ? io_r_109_b : _GEN_18688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18690 = 9'h6e == r_count_46_io_out ? io_r_110_b : _GEN_18689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18691 = 9'h6f == r_count_46_io_out ? io_r_111_b : _GEN_18690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18692 = 9'h70 == r_count_46_io_out ? io_r_112_b : _GEN_18691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18693 = 9'h71 == r_count_46_io_out ? io_r_113_b : _GEN_18692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18694 = 9'h72 == r_count_46_io_out ? io_r_114_b : _GEN_18693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18695 = 9'h73 == r_count_46_io_out ? io_r_115_b : _GEN_18694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18696 = 9'h74 == r_count_46_io_out ? io_r_116_b : _GEN_18695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18697 = 9'h75 == r_count_46_io_out ? io_r_117_b : _GEN_18696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18698 = 9'h76 == r_count_46_io_out ? io_r_118_b : _GEN_18697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18699 = 9'h77 == r_count_46_io_out ? io_r_119_b : _GEN_18698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18700 = 9'h78 == r_count_46_io_out ? io_r_120_b : _GEN_18699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18701 = 9'h79 == r_count_46_io_out ? io_r_121_b : _GEN_18700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18702 = 9'h7a == r_count_46_io_out ? io_r_122_b : _GEN_18701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18703 = 9'h7b == r_count_46_io_out ? io_r_123_b : _GEN_18702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18704 = 9'h7c == r_count_46_io_out ? io_r_124_b : _GEN_18703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18705 = 9'h7d == r_count_46_io_out ? io_r_125_b : _GEN_18704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18706 = 9'h7e == r_count_46_io_out ? io_r_126_b : _GEN_18705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18707 = 9'h7f == r_count_46_io_out ? io_r_127_b : _GEN_18706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18708 = 9'h80 == r_count_46_io_out ? io_r_128_b : _GEN_18707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18709 = 9'h81 == r_count_46_io_out ? io_r_129_b : _GEN_18708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18710 = 9'h82 == r_count_46_io_out ? io_r_130_b : _GEN_18709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18711 = 9'h83 == r_count_46_io_out ? io_r_131_b : _GEN_18710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18712 = 9'h84 == r_count_46_io_out ? io_r_132_b : _GEN_18711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18713 = 9'h85 == r_count_46_io_out ? io_r_133_b : _GEN_18712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18714 = 9'h86 == r_count_46_io_out ? io_r_134_b : _GEN_18713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18715 = 9'h87 == r_count_46_io_out ? io_r_135_b : _GEN_18714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18716 = 9'h88 == r_count_46_io_out ? io_r_136_b : _GEN_18715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18717 = 9'h89 == r_count_46_io_out ? io_r_137_b : _GEN_18716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18718 = 9'h8a == r_count_46_io_out ? io_r_138_b : _GEN_18717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18719 = 9'h8b == r_count_46_io_out ? io_r_139_b : _GEN_18718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18720 = 9'h8c == r_count_46_io_out ? io_r_140_b : _GEN_18719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18721 = 9'h8d == r_count_46_io_out ? io_r_141_b : _GEN_18720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18722 = 9'h8e == r_count_46_io_out ? io_r_142_b : _GEN_18721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18723 = 9'h8f == r_count_46_io_out ? io_r_143_b : _GEN_18722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18724 = 9'h90 == r_count_46_io_out ? io_r_144_b : _GEN_18723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18725 = 9'h91 == r_count_46_io_out ? io_r_145_b : _GEN_18724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18726 = 9'h92 == r_count_46_io_out ? io_r_146_b : _GEN_18725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18727 = 9'h93 == r_count_46_io_out ? io_r_147_b : _GEN_18726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18728 = 9'h94 == r_count_46_io_out ? io_r_148_b : _GEN_18727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18729 = 9'h95 == r_count_46_io_out ? io_r_149_b : _GEN_18728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18730 = 9'h96 == r_count_46_io_out ? io_r_150_b : _GEN_18729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18731 = 9'h97 == r_count_46_io_out ? io_r_151_b : _GEN_18730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18732 = 9'h98 == r_count_46_io_out ? io_r_152_b : _GEN_18731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18733 = 9'h99 == r_count_46_io_out ? io_r_153_b : _GEN_18732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18734 = 9'h9a == r_count_46_io_out ? io_r_154_b : _GEN_18733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18735 = 9'h9b == r_count_46_io_out ? io_r_155_b : _GEN_18734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18736 = 9'h9c == r_count_46_io_out ? io_r_156_b : _GEN_18735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18737 = 9'h9d == r_count_46_io_out ? io_r_157_b : _GEN_18736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18738 = 9'h9e == r_count_46_io_out ? io_r_158_b : _GEN_18737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18739 = 9'h9f == r_count_46_io_out ? io_r_159_b : _GEN_18738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18740 = 9'ha0 == r_count_46_io_out ? io_r_160_b : _GEN_18739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18741 = 9'ha1 == r_count_46_io_out ? io_r_161_b : _GEN_18740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18742 = 9'ha2 == r_count_46_io_out ? io_r_162_b : _GEN_18741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18743 = 9'ha3 == r_count_46_io_out ? io_r_163_b : _GEN_18742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18744 = 9'ha4 == r_count_46_io_out ? io_r_164_b : _GEN_18743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18745 = 9'ha5 == r_count_46_io_out ? io_r_165_b : _GEN_18744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18746 = 9'ha6 == r_count_46_io_out ? io_r_166_b : _GEN_18745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18747 = 9'ha7 == r_count_46_io_out ? io_r_167_b : _GEN_18746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18748 = 9'ha8 == r_count_46_io_out ? io_r_168_b : _GEN_18747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18749 = 9'ha9 == r_count_46_io_out ? io_r_169_b : _GEN_18748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18750 = 9'haa == r_count_46_io_out ? io_r_170_b : _GEN_18749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18751 = 9'hab == r_count_46_io_out ? io_r_171_b : _GEN_18750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18752 = 9'hac == r_count_46_io_out ? io_r_172_b : _GEN_18751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18753 = 9'had == r_count_46_io_out ? io_r_173_b : _GEN_18752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18754 = 9'hae == r_count_46_io_out ? io_r_174_b : _GEN_18753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18755 = 9'haf == r_count_46_io_out ? io_r_175_b : _GEN_18754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18756 = 9'hb0 == r_count_46_io_out ? io_r_176_b : _GEN_18755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18757 = 9'hb1 == r_count_46_io_out ? io_r_177_b : _GEN_18756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18758 = 9'hb2 == r_count_46_io_out ? io_r_178_b : _GEN_18757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18759 = 9'hb3 == r_count_46_io_out ? io_r_179_b : _GEN_18758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18760 = 9'hb4 == r_count_46_io_out ? io_r_180_b : _GEN_18759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18761 = 9'hb5 == r_count_46_io_out ? io_r_181_b : _GEN_18760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18762 = 9'hb6 == r_count_46_io_out ? io_r_182_b : _GEN_18761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18763 = 9'hb7 == r_count_46_io_out ? io_r_183_b : _GEN_18762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18764 = 9'hb8 == r_count_46_io_out ? io_r_184_b : _GEN_18763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18765 = 9'hb9 == r_count_46_io_out ? io_r_185_b : _GEN_18764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18766 = 9'hba == r_count_46_io_out ? io_r_186_b : _GEN_18765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18767 = 9'hbb == r_count_46_io_out ? io_r_187_b : _GEN_18766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18768 = 9'hbc == r_count_46_io_out ? io_r_188_b : _GEN_18767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18769 = 9'hbd == r_count_46_io_out ? io_r_189_b : _GEN_18768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18770 = 9'hbe == r_count_46_io_out ? io_r_190_b : _GEN_18769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18771 = 9'hbf == r_count_46_io_out ? io_r_191_b : _GEN_18770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18772 = 9'hc0 == r_count_46_io_out ? io_r_192_b : _GEN_18771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18773 = 9'hc1 == r_count_46_io_out ? io_r_193_b : _GEN_18772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18774 = 9'hc2 == r_count_46_io_out ? io_r_194_b : _GEN_18773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18775 = 9'hc3 == r_count_46_io_out ? io_r_195_b : _GEN_18774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18776 = 9'hc4 == r_count_46_io_out ? io_r_196_b : _GEN_18775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18777 = 9'hc5 == r_count_46_io_out ? io_r_197_b : _GEN_18776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18778 = 9'hc6 == r_count_46_io_out ? io_r_198_b : _GEN_18777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18779 = 9'hc7 == r_count_46_io_out ? io_r_199_b : _GEN_18778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18780 = 9'hc8 == r_count_46_io_out ? io_r_200_b : _GEN_18779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18781 = 9'hc9 == r_count_46_io_out ? io_r_201_b : _GEN_18780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18782 = 9'hca == r_count_46_io_out ? io_r_202_b : _GEN_18781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18783 = 9'hcb == r_count_46_io_out ? io_r_203_b : _GEN_18782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18784 = 9'hcc == r_count_46_io_out ? io_r_204_b : _GEN_18783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18785 = 9'hcd == r_count_46_io_out ? io_r_205_b : _GEN_18784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18786 = 9'hce == r_count_46_io_out ? io_r_206_b : _GEN_18785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18787 = 9'hcf == r_count_46_io_out ? io_r_207_b : _GEN_18786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18788 = 9'hd0 == r_count_46_io_out ? io_r_208_b : _GEN_18787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18789 = 9'hd1 == r_count_46_io_out ? io_r_209_b : _GEN_18788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18790 = 9'hd2 == r_count_46_io_out ? io_r_210_b : _GEN_18789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18791 = 9'hd3 == r_count_46_io_out ? io_r_211_b : _GEN_18790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18792 = 9'hd4 == r_count_46_io_out ? io_r_212_b : _GEN_18791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18793 = 9'hd5 == r_count_46_io_out ? io_r_213_b : _GEN_18792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18794 = 9'hd6 == r_count_46_io_out ? io_r_214_b : _GEN_18793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18795 = 9'hd7 == r_count_46_io_out ? io_r_215_b : _GEN_18794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18796 = 9'hd8 == r_count_46_io_out ? io_r_216_b : _GEN_18795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18797 = 9'hd9 == r_count_46_io_out ? io_r_217_b : _GEN_18796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18798 = 9'hda == r_count_46_io_out ? io_r_218_b : _GEN_18797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18799 = 9'hdb == r_count_46_io_out ? io_r_219_b : _GEN_18798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18800 = 9'hdc == r_count_46_io_out ? io_r_220_b : _GEN_18799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18801 = 9'hdd == r_count_46_io_out ? io_r_221_b : _GEN_18800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18802 = 9'hde == r_count_46_io_out ? io_r_222_b : _GEN_18801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18803 = 9'hdf == r_count_46_io_out ? io_r_223_b : _GEN_18802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18804 = 9'he0 == r_count_46_io_out ? io_r_224_b : _GEN_18803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18805 = 9'he1 == r_count_46_io_out ? io_r_225_b : _GEN_18804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18806 = 9'he2 == r_count_46_io_out ? io_r_226_b : _GEN_18805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18807 = 9'he3 == r_count_46_io_out ? io_r_227_b : _GEN_18806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18808 = 9'he4 == r_count_46_io_out ? io_r_228_b : _GEN_18807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18809 = 9'he5 == r_count_46_io_out ? io_r_229_b : _GEN_18808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18810 = 9'he6 == r_count_46_io_out ? io_r_230_b : _GEN_18809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18811 = 9'he7 == r_count_46_io_out ? io_r_231_b : _GEN_18810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18812 = 9'he8 == r_count_46_io_out ? io_r_232_b : _GEN_18811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18813 = 9'he9 == r_count_46_io_out ? io_r_233_b : _GEN_18812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18814 = 9'hea == r_count_46_io_out ? io_r_234_b : _GEN_18813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18815 = 9'heb == r_count_46_io_out ? io_r_235_b : _GEN_18814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18816 = 9'hec == r_count_46_io_out ? io_r_236_b : _GEN_18815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18817 = 9'hed == r_count_46_io_out ? io_r_237_b : _GEN_18816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18818 = 9'hee == r_count_46_io_out ? io_r_238_b : _GEN_18817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18819 = 9'hef == r_count_46_io_out ? io_r_239_b : _GEN_18818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18820 = 9'hf0 == r_count_46_io_out ? io_r_240_b : _GEN_18819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18821 = 9'hf1 == r_count_46_io_out ? io_r_241_b : _GEN_18820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18822 = 9'hf2 == r_count_46_io_out ? io_r_242_b : _GEN_18821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18823 = 9'hf3 == r_count_46_io_out ? io_r_243_b : _GEN_18822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18824 = 9'hf4 == r_count_46_io_out ? io_r_244_b : _GEN_18823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18825 = 9'hf5 == r_count_46_io_out ? io_r_245_b : _GEN_18824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18826 = 9'hf6 == r_count_46_io_out ? io_r_246_b : _GEN_18825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18827 = 9'hf7 == r_count_46_io_out ? io_r_247_b : _GEN_18826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18828 = 9'hf8 == r_count_46_io_out ? io_r_248_b : _GEN_18827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18829 = 9'hf9 == r_count_46_io_out ? io_r_249_b : _GEN_18828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18830 = 9'hfa == r_count_46_io_out ? io_r_250_b : _GEN_18829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18831 = 9'hfb == r_count_46_io_out ? io_r_251_b : _GEN_18830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18832 = 9'hfc == r_count_46_io_out ? io_r_252_b : _GEN_18831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18833 = 9'hfd == r_count_46_io_out ? io_r_253_b : _GEN_18832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18834 = 9'hfe == r_count_46_io_out ? io_r_254_b : _GEN_18833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18835 = 9'hff == r_count_46_io_out ? io_r_255_b : _GEN_18834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18836 = 9'h100 == r_count_46_io_out ? io_r_256_b : _GEN_18835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18837 = 9'h101 == r_count_46_io_out ? io_r_257_b : _GEN_18836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18838 = 9'h102 == r_count_46_io_out ? io_r_258_b : _GEN_18837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18839 = 9'h103 == r_count_46_io_out ? io_r_259_b : _GEN_18838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18840 = 9'h104 == r_count_46_io_out ? io_r_260_b : _GEN_18839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18841 = 9'h105 == r_count_46_io_out ? io_r_261_b : _GEN_18840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18842 = 9'h106 == r_count_46_io_out ? io_r_262_b : _GEN_18841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18843 = 9'h107 == r_count_46_io_out ? io_r_263_b : _GEN_18842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18844 = 9'h108 == r_count_46_io_out ? io_r_264_b : _GEN_18843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18845 = 9'h109 == r_count_46_io_out ? io_r_265_b : _GEN_18844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18846 = 9'h10a == r_count_46_io_out ? io_r_266_b : _GEN_18845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18847 = 9'h10b == r_count_46_io_out ? io_r_267_b : _GEN_18846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18848 = 9'h10c == r_count_46_io_out ? io_r_268_b : _GEN_18847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18849 = 9'h10d == r_count_46_io_out ? io_r_269_b : _GEN_18848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18850 = 9'h10e == r_count_46_io_out ? io_r_270_b : _GEN_18849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18851 = 9'h10f == r_count_46_io_out ? io_r_271_b : _GEN_18850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18852 = 9'h110 == r_count_46_io_out ? io_r_272_b : _GEN_18851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18853 = 9'h111 == r_count_46_io_out ? io_r_273_b : _GEN_18852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18854 = 9'h112 == r_count_46_io_out ? io_r_274_b : _GEN_18853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18855 = 9'h113 == r_count_46_io_out ? io_r_275_b : _GEN_18854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18856 = 9'h114 == r_count_46_io_out ? io_r_276_b : _GEN_18855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18857 = 9'h115 == r_count_46_io_out ? io_r_277_b : _GEN_18856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18858 = 9'h116 == r_count_46_io_out ? io_r_278_b : _GEN_18857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18859 = 9'h117 == r_count_46_io_out ? io_r_279_b : _GEN_18858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18860 = 9'h118 == r_count_46_io_out ? io_r_280_b : _GEN_18859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18861 = 9'h119 == r_count_46_io_out ? io_r_281_b : _GEN_18860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18862 = 9'h11a == r_count_46_io_out ? io_r_282_b : _GEN_18861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18863 = 9'h11b == r_count_46_io_out ? io_r_283_b : _GEN_18862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18864 = 9'h11c == r_count_46_io_out ? io_r_284_b : _GEN_18863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18865 = 9'h11d == r_count_46_io_out ? io_r_285_b : _GEN_18864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18866 = 9'h11e == r_count_46_io_out ? io_r_286_b : _GEN_18865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18867 = 9'h11f == r_count_46_io_out ? io_r_287_b : _GEN_18866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18868 = 9'h120 == r_count_46_io_out ? io_r_288_b : _GEN_18867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18869 = 9'h121 == r_count_46_io_out ? io_r_289_b : _GEN_18868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18870 = 9'h122 == r_count_46_io_out ? io_r_290_b : _GEN_18869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18871 = 9'h123 == r_count_46_io_out ? io_r_291_b : _GEN_18870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18872 = 9'h124 == r_count_46_io_out ? io_r_292_b : _GEN_18871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18873 = 9'h125 == r_count_46_io_out ? io_r_293_b : _GEN_18872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18874 = 9'h126 == r_count_46_io_out ? io_r_294_b : _GEN_18873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18875 = 9'h127 == r_count_46_io_out ? io_r_295_b : _GEN_18874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18876 = 9'h128 == r_count_46_io_out ? io_r_296_b : _GEN_18875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18877 = 9'h129 == r_count_46_io_out ? io_r_297_b : _GEN_18876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18878 = 9'h12a == r_count_46_io_out ? io_r_298_b : _GEN_18877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18879 = 9'h12b == r_count_46_io_out ? io_r_299_b : _GEN_18878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18880 = 9'h12c == r_count_46_io_out ? io_r_300_b : _GEN_18879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18881 = 9'h12d == r_count_46_io_out ? io_r_301_b : _GEN_18880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18882 = 9'h12e == r_count_46_io_out ? io_r_302_b : _GEN_18881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18883 = 9'h12f == r_count_46_io_out ? io_r_303_b : _GEN_18882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18884 = 9'h130 == r_count_46_io_out ? io_r_304_b : _GEN_18883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18885 = 9'h131 == r_count_46_io_out ? io_r_305_b : _GEN_18884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18886 = 9'h132 == r_count_46_io_out ? io_r_306_b : _GEN_18885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18887 = 9'h133 == r_count_46_io_out ? io_r_307_b : _GEN_18886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18888 = 9'h134 == r_count_46_io_out ? io_r_308_b : _GEN_18887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18889 = 9'h135 == r_count_46_io_out ? io_r_309_b : _GEN_18888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18890 = 9'h136 == r_count_46_io_out ? io_r_310_b : _GEN_18889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18891 = 9'h137 == r_count_46_io_out ? io_r_311_b : _GEN_18890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18892 = 9'h138 == r_count_46_io_out ? io_r_312_b : _GEN_18891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18893 = 9'h139 == r_count_46_io_out ? io_r_313_b : _GEN_18892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18894 = 9'h13a == r_count_46_io_out ? io_r_314_b : _GEN_18893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18895 = 9'h13b == r_count_46_io_out ? io_r_315_b : _GEN_18894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18896 = 9'h13c == r_count_46_io_out ? io_r_316_b : _GEN_18895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18897 = 9'h13d == r_count_46_io_out ? io_r_317_b : _GEN_18896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18898 = 9'h13e == r_count_46_io_out ? io_r_318_b : _GEN_18897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18899 = 9'h13f == r_count_46_io_out ? io_r_319_b : _GEN_18898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18900 = 9'h140 == r_count_46_io_out ? io_r_320_b : _GEN_18899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18901 = 9'h141 == r_count_46_io_out ? io_r_321_b : _GEN_18900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18902 = 9'h142 == r_count_46_io_out ? io_r_322_b : _GEN_18901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18903 = 9'h143 == r_count_46_io_out ? io_r_323_b : _GEN_18902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18904 = 9'h144 == r_count_46_io_out ? io_r_324_b : _GEN_18903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18905 = 9'h145 == r_count_46_io_out ? io_r_325_b : _GEN_18904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18906 = 9'h146 == r_count_46_io_out ? io_r_326_b : _GEN_18905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18907 = 9'h147 == r_count_46_io_out ? io_r_327_b : _GEN_18906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18908 = 9'h148 == r_count_46_io_out ? io_r_328_b : _GEN_18907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18909 = 9'h149 == r_count_46_io_out ? io_r_329_b : _GEN_18908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18910 = 9'h14a == r_count_46_io_out ? io_r_330_b : _GEN_18909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18911 = 9'h14b == r_count_46_io_out ? io_r_331_b : _GEN_18910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18912 = 9'h14c == r_count_46_io_out ? io_r_332_b : _GEN_18911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18913 = 9'h14d == r_count_46_io_out ? io_r_333_b : _GEN_18912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18914 = 9'h14e == r_count_46_io_out ? io_r_334_b : _GEN_18913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18915 = 9'h14f == r_count_46_io_out ? io_r_335_b : _GEN_18914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18916 = 9'h150 == r_count_46_io_out ? io_r_336_b : _GEN_18915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18917 = 9'h151 == r_count_46_io_out ? io_r_337_b : _GEN_18916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18918 = 9'h152 == r_count_46_io_out ? io_r_338_b : _GEN_18917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18919 = 9'h153 == r_count_46_io_out ? io_r_339_b : _GEN_18918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18920 = 9'h154 == r_count_46_io_out ? io_r_340_b : _GEN_18919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18921 = 9'h155 == r_count_46_io_out ? io_r_341_b : _GEN_18920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18922 = 9'h156 == r_count_46_io_out ? io_r_342_b : _GEN_18921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18923 = 9'h157 == r_count_46_io_out ? io_r_343_b : _GEN_18922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18924 = 9'h158 == r_count_46_io_out ? io_r_344_b : _GEN_18923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18925 = 9'h159 == r_count_46_io_out ? io_r_345_b : _GEN_18924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18926 = 9'h15a == r_count_46_io_out ? io_r_346_b : _GEN_18925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18927 = 9'h15b == r_count_46_io_out ? io_r_347_b : _GEN_18926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18928 = 9'h15c == r_count_46_io_out ? io_r_348_b : _GEN_18927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18929 = 9'h15d == r_count_46_io_out ? io_r_349_b : _GEN_18928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18930 = 9'h15e == r_count_46_io_out ? io_r_350_b : _GEN_18929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18931 = 9'h15f == r_count_46_io_out ? io_r_351_b : _GEN_18930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18932 = 9'h160 == r_count_46_io_out ? io_r_352_b : _GEN_18931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18933 = 9'h161 == r_count_46_io_out ? io_r_353_b : _GEN_18932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18934 = 9'h162 == r_count_46_io_out ? io_r_354_b : _GEN_18933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18935 = 9'h163 == r_count_46_io_out ? io_r_355_b : _GEN_18934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18936 = 9'h164 == r_count_46_io_out ? io_r_356_b : _GEN_18935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18937 = 9'h165 == r_count_46_io_out ? io_r_357_b : _GEN_18936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18938 = 9'h166 == r_count_46_io_out ? io_r_358_b : _GEN_18937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18939 = 9'h167 == r_count_46_io_out ? io_r_359_b : _GEN_18938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18940 = 9'h168 == r_count_46_io_out ? io_r_360_b : _GEN_18939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18941 = 9'h169 == r_count_46_io_out ? io_r_361_b : _GEN_18940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18942 = 9'h16a == r_count_46_io_out ? io_r_362_b : _GEN_18941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18943 = 9'h16b == r_count_46_io_out ? io_r_363_b : _GEN_18942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18944 = 9'h16c == r_count_46_io_out ? io_r_364_b : _GEN_18943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18945 = 9'h16d == r_count_46_io_out ? io_r_365_b : _GEN_18944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18946 = 9'h16e == r_count_46_io_out ? io_r_366_b : _GEN_18945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18947 = 9'h16f == r_count_46_io_out ? io_r_367_b : _GEN_18946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18948 = 9'h170 == r_count_46_io_out ? io_r_368_b : _GEN_18947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18949 = 9'h171 == r_count_46_io_out ? io_r_369_b : _GEN_18948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18950 = 9'h172 == r_count_46_io_out ? io_r_370_b : _GEN_18949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18951 = 9'h173 == r_count_46_io_out ? io_r_371_b : _GEN_18950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18952 = 9'h174 == r_count_46_io_out ? io_r_372_b : _GEN_18951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18953 = 9'h175 == r_count_46_io_out ? io_r_373_b : _GEN_18952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18954 = 9'h176 == r_count_46_io_out ? io_r_374_b : _GEN_18953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18955 = 9'h177 == r_count_46_io_out ? io_r_375_b : _GEN_18954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18956 = 9'h178 == r_count_46_io_out ? io_r_376_b : _GEN_18955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18957 = 9'h179 == r_count_46_io_out ? io_r_377_b : _GEN_18956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18958 = 9'h17a == r_count_46_io_out ? io_r_378_b : _GEN_18957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18959 = 9'h17b == r_count_46_io_out ? io_r_379_b : _GEN_18958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18960 = 9'h17c == r_count_46_io_out ? io_r_380_b : _GEN_18959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18961 = 9'h17d == r_count_46_io_out ? io_r_381_b : _GEN_18960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18962 = 9'h17e == r_count_46_io_out ? io_r_382_b : _GEN_18961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18963 = 9'h17f == r_count_46_io_out ? io_r_383_b : _GEN_18962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18964 = 9'h180 == r_count_46_io_out ? io_r_384_b : _GEN_18963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18965 = 9'h181 == r_count_46_io_out ? io_r_385_b : _GEN_18964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18966 = 9'h182 == r_count_46_io_out ? io_r_386_b : _GEN_18965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18967 = 9'h183 == r_count_46_io_out ? io_r_387_b : _GEN_18966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18968 = 9'h184 == r_count_46_io_out ? io_r_388_b : _GEN_18967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18969 = 9'h185 == r_count_46_io_out ? io_r_389_b : _GEN_18968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18970 = 9'h186 == r_count_46_io_out ? io_r_390_b : _GEN_18969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18971 = 9'h187 == r_count_46_io_out ? io_r_391_b : _GEN_18970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18972 = 9'h188 == r_count_46_io_out ? io_r_392_b : _GEN_18971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18973 = 9'h189 == r_count_46_io_out ? io_r_393_b : _GEN_18972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18974 = 9'h18a == r_count_46_io_out ? io_r_394_b : _GEN_18973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18975 = 9'h18b == r_count_46_io_out ? io_r_395_b : _GEN_18974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18976 = 9'h18c == r_count_46_io_out ? io_r_396_b : _GEN_18975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18977 = 9'h18d == r_count_46_io_out ? io_r_397_b : _GEN_18976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18978 = 9'h18e == r_count_46_io_out ? io_r_398_b : _GEN_18977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18981 = 9'h1 == r_count_47_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18982 = 9'h2 == r_count_47_io_out ? io_r_2_b : _GEN_18981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18983 = 9'h3 == r_count_47_io_out ? io_r_3_b : _GEN_18982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18984 = 9'h4 == r_count_47_io_out ? io_r_4_b : _GEN_18983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18985 = 9'h5 == r_count_47_io_out ? io_r_5_b : _GEN_18984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18986 = 9'h6 == r_count_47_io_out ? io_r_6_b : _GEN_18985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18987 = 9'h7 == r_count_47_io_out ? io_r_7_b : _GEN_18986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18988 = 9'h8 == r_count_47_io_out ? io_r_8_b : _GEN_18987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18989 = 9'h9 == r_count_47_io_out ? io_r_9_b : _GEN_18988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18990 = 9'ha == r_count_47_io_out ? io_r_10_b : _GEN_18989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18991 = 9'hb == r_count_47_io_out ? io_r_11_b : _GEN_18990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18992 = 9'hc == r_count_47_io_out ? io_r_12_b : _GEN_18991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18993 = 9'hd == r_count_47_io_out ? io_r_13_b : _GEN_18992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18994 = 9'he == r_count_47_io_out ? io_r_14_b : _GEN_18993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18995 = 9'hf == r_count_47_io_out ? io_r_15_b : _GEN_18994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18996 = 9'h10 == r_count_47_io_out ? io_r_16_b : _GEN_18995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18997 = 9'h11 == r_count_47_io_out ? io_r_17_b : _GEN_18996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18998 = 9'h12 == r_count_47_io_out ? io_r_18_b : _GEN_18997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18999 = 9'h13 == r_count_47_io_out ? io_r_19_b : _GEN_18998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19000 = 9'h14 == r_count_47_io_out ? io_r_20_b : _GEN_18999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19001 = 9'h15 == r_count_47_io_out ? io_r_21_b : _GEN_19000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19002 = 9'h16 == r_count_47_io_out ? io_r_22_b : _GEN_19001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19003 = 9'h17 == r_count_47_io_out ? io_r_23_b : _GEN_19002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19004 = 9'h18 == r_count_47_io_out ? io_r_24_b : _GEN_19003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19005 = 9'h19 == r_count_47_io_out ? io_r_25_b : _GEN_19004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19006 = 9'h1a == r_count_47_io_out ? io_r_26_b : _GEN_19005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19007 = 9'h1b == r_count_47_io_out ? io_r_27_b : _GEN_19006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19008 = 9'h1c == r_count_47_io_out ? io_r_28_b : _GEN_19007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19009 = 9'h1d == r_count_47_io_out ? io_r_29_b : _GEN_19008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19010 = 9'h1e == r_count_47_io_out ? io_r_30_b : _GEN_19009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19011 = 9'h1f == r_count_47_io_out ? io_r_31_b : _GEN_19010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19012 = 9'h20 == r_count_47_io_out ? io_r_32_b : _GEN_19011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19013 = 9'h21 == r_count_47_io_out ? io_r_33_b : _GEN_19012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19014 = 9'h22 == r_count_47_io_out ? io_r_34_b : _GEN_19013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19015 = 9'h23 == r_count_47_io_out ? io_r_35_b : _GEN_19014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19016 = 9'h24 == r_count_47_io_out ? io_r_36_b : _GEN_19015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19017 = 9'h25 == r_count_47_io_out ? io_r_37_b : _GEN_19016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19018 = 9'h26 == r_count_47_io_out ? io_r_38_b : _GEN_19017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19019 = 9'h27 == r_count_47_io_out ? io_r_39_b : _GEN_19018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19020 = 9'h28 == r_count_47_io_out ? io_r_40_b : _GEN_19019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19021 = 9'h29 == r_count_47_io_out ? io_r_41_b : _GEN_19020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19022 = 9'h2a == r_count_47_io_out ? io_r_42_b : _GEN_19021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19023 = 9'h2b == r_count_47_io_out ? io_r_43_b : _GEN_19022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19024 = 9'h2c == r_count_47_io_out ? io_r_44_b : _GEN_19023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19025 = 9'h2d == r_count_47_io_out ? io_r_45_b : _GEN_19024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19026 = 9'h2e == r_count_47_io_out ? io_r_46_b : _GEN_19025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19027 = 9'h2f == r_count_47_io_out ? io_r_47_b : _GEN_19026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19028 = 9'h30 == r_count_47_io_out ? io_r_48_b : _GEN_19027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19029 = 9'h31 == r_count_47_io_out ? io_r_49_b : _GEN_19028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19030 = 9'h32 == r_count_47_io_out ? io_r_50_b : _GEN_19029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19031 = 9'h33 == r_count_47_io_out ? io_r_51_b : _GEN_19030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19032 = 9'h34 == r_count_47_io_out ? io_r_52_b : _GEN_19031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19033 = 9'h35 == r_count_47_io_out ? io_r_53_b : _GEN_19032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19034 = 9'h36 == r_count_47_io_out ? io_r_54_b : _GEN_19033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19035 = 9'h37 == r_count_47_io_out ? io_r_55_b : _GEN_19034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19036 = 9'h38 == r_count_47_io_out ? io_r_56_b : _GEN_19035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19037 = 9'h39 == r_count_47_io_out ? io_r_57_b : _GEN_19036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19038 = 9'h3a == r_count_47_io_out ? io_r_58_b : _GEN_19037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19039 = 9'h3b == r_count_47_io_out ? io_r_59_b : _GEN_19038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19040 = 9'h3c == r_count_47_io_out ? io_r_60_b : _GEN_19039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19041 = 9'h3d == r_count_47_io_out ? io_r_61_b : _GEN_19040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19042 = 9'h3e == r_count_47_io_out ? io_r_62_b : _GEN_19041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19043 = 9'h3f == r_count_47_io_out ? io_r_63_b : _GEN_19042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19044 = 9'h40 == r_count_47_io_out ? io_r_64_b : _GEN_19043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19045 = 9'h41 == r_count_47_io_out ? io_r_65_b : _GEN_19044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19046 = 9'h42 == r_count_47_io_out ? io_r_66_b : _GEN_19045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19047 = 9'h43 == r_count_47_io_out ? io_r_67_b : _GEN_19046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19048 = 9'h44 == r_count_47_io_out ? io_r_68_b : _GEN_19047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19049 = 9'h45 == r_count_47_io_out ? io_r_69_b : _GEN_19048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19050 = 9'h46 == r_count_47_io_out ? io_r_70_b : _GEN_19049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19051 = 9'h47 == r_count_47_io_out ? io_r_71_b : _GEN_19050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19052 = 9'h48 == r_count_47_io_out ? io_r_72_b : _GEN_19051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19053 = 9'h49 == r_count_47_io_out ? io_r_73_b : _GEN_19052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19054 = 9'h4a == r_count_47_io_out ? io_r_74_b : _GEN_19053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19055 = 9'h4b == r_count_47_io_out ? io_r_75_b : _GEN_19054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19056 = 9'h4c == r_count_47_io_out ? io_r_76_b : _GEN_19055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19057 = 9'h4d == r_count_47_io_out ? io_r_77_b : _GEN_19056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19058 = 9'h4e == r_count_47_io_out ? io_r_78_b : _GEN_19057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19059 = 9'h4f == r_count_47_io_out ? io_r_79_b : _GEN_19058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19060 = 9'h50 == r_count_47_io_out ? io_r_80_b : _GEN_19059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19061 = 9'h51 == r_count_47_io_out ? io_r_81_b : _GEN_19060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19062 = 9'h52 == r_count_47_io_out ? io_r_82_b : _GEN_19061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19063 = 9'h53 == r_count_47_io_out ? io_r_83_b : _GEN_19062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19064 = 9'h54 == r_count_47_io_out ? io_r_84_b : _GEN_19063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19065 = 9'h55 == r_count_47_io_out ? io_r_85_b : _GEN_19064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19066 = 9'h56 == r_count_47_io_out ? io_r_86_b : _GEN_19065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19067 = 9'h57 == r_count_47_io_out ? io_r_87_b : _GEN_19066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19068 = 9'h58 == r_count_47_io_out ? io_r_88_b : _GEN_19067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19069 = 9'h59 == r_count_47_io_out ? io_r_89_b : _GEN_19068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19070 = 9'h5a == r_count_47_io_out ? io_r_90_b : _GEN_19069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19071 = 9'h5b == r_count_47_io_out ? io_r_91_b : _GEN_19070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19072 = 9'h5c == r_count_47_io_out ? io_r_92_b : _GEN_19071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19073 = 9'h5d == r_count_47_io_out ? io_r_93_b : _GEN_19072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19074 = 9'h5e == r_count_47_io_out ? io_r_94_b : _GEN_19073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19075 = 9'h5f == r_count_47_io_out ? io_r_95_b : _GEN_19074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19076 = 9'h60 == r_count_47_io_out ? io_r_96_b : _GEN_19075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19077 = 9'h61 == r_count_47_io_out ? io_r_97_b : _GEN_19076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19078 = 9'h62 == r_count_47_io_out ? io_r_98_b : _GEN_19077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19079 = 9'h63 == r_count_47_io_out ? io_r_99_b : _GEN_19078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19080 = 9'h64 == r_count_47_io_out ? io_r_100_b : _GEN_19079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19081 = 9'h65 == r_count_47_io_out ? io_r_101_b : _GEN_19080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19082 = 9'h66 == r_count_47_io_out ? io_r_102_b : _GEN_19081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19083 = 9'h67 == r_count_47_io_out ? io_r_103_b : _GEN_19082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19084 = 9'h68 == r_count_47_io_out ? io_r_104_b : _GEN_19083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19085 = 9'h69 == r_count_47_io_out ? io_r_105_b : _GEN_19084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19086 = 9'h6a == r_count_47_io_out ? io_r_106_b : _GEN_19085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19087 = 9'h6b == r_count_47_io_out ? io_r_107_b : _GEN_19086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19088 = 9'h6c == r_count_47_io_out ? io_r_108_b : _GEN_19087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19089 = 9'h6d == r_count_47_io_out ? io_r_109_b : _GEN_19088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19090 = 9'h6e == r_count_47_io_out ? io_r_110_b : _GEN_19089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19091 = 9'h6f == r_count_47_io_out ? io_r_111_b : _GEN_19090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19092 = 9'h70 == r_count_47_io_out ? io_r_112_b : _GEN_19091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19093 = 9'h71 == r_count_47_io_out ? io_r_113_b : _GEN_19092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19094 = 9'h72 == r_count_47_io_out ? io_r_114_b : _GEN_19093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19095 = 9'h73 == r_count_47_io_out ? io_r_115_b : _GEN_19094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19096 = 9'h74 == r_count_47_io_out ? io_r_116_b : _GEN_19095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19097 = 9'h75 == r_count_47_io_out ? io_r_117_b : _GEN_19096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19098 = 9'h76 == r_count_47_io_out ? io_r_118_b : _GEN_19097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19099 = 9'h77 == r_count_47_io_out ? io_r_119_b : _GEN_19098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19100 = 9'h78 == r_count_47_io_out ? io_r_120_b : _GEN_19099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19101 = 9'h79 == r_count_47_io_out ? io_r_121_b : _GEN_19100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19102 = 9'h7a == r_count_47_io_out ? io_r_122_b : _GEN_19101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19103 = 9'h7b == r_count_47_io_out ? io_r_123_b : _GEN_19102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19104 = 9'h7c == r_count_47_io_out ? io_r_124_b : _GEN_19103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19105 = 9'h7d == r_count_47_io_out ? io_r_125_b : _GEN_19104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19106 = 9'h7e == r_count_47_io_out ? io_r_126_b : _GEN_19105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19107 = 9'h7f == r_count_47_io_out ? io_r_127_b : _GEN_19106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19108 = 9'h80 == r_count_47_io_out ? io_r_128_b : _GEN_19107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19109 = 9'h81 == r_count_47_io_out ? io_r_129_b : _GEN_19108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19110 = 9'h82 == r_count_47_io_out ? io_r_130_b : _GEN_19109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19111 = 9'h83 == r_count_47_io_out ? io_r_131_b : _GEN_19110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19112 = 9'h84 == r_count_47_io_out ? io_r_132_b : _GEN_19111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19113 = 9'h85 == r_count_47_io_out ? io_r_133_b : _GEN_19112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19114 = 9'h86 == r_count_47_io_out ? io_r_134_b : _GEN_19113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19115 = 9'h87 == r_count_47_io_out ? io_r_135_b : _GEN_19114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19116 = 9'h88 == r_count_47_io_out ? io_r_136_b : _GEN_19115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19117 = 9'h89 == r_count_47_io_out ? io_r_137_b : _GEN_19116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19118 = 9'h8a == r_count_47_io_out ? io_r_138_b : _GEN_19117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19119 = 9'h8b == r_count_47_io_out ? io_r_139_b : _GEN_19118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19120 = 9'h8c == r_count_47_io_out ? io_r_140_b : _GEN_19119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19121 = 9'h8d == r_count_47_io_out ? io_r_141_b : _GEN_19120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19122 = 9'h8e == r_count_47_io_out ? io_r_142_b : _GEN_19121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19123 = 9'h8f == r_count_47_io_out ? io_r_143_b : _GEN_19122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19124 = 9'h90 == r_count_47_io_out ? io_r_144_b : _GEN_19123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19125 = 9'h91 == r_count_47_io_out ? io_r_145_b : _GEN_19124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19126 = 9'h92 == r_count_47_io_out ? io_r_146_b : _GEN_19125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19127 = 9'h93 == r_count_47_io_out ? io_r_147_b : _GEN_19126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19128 = 9'h94 == r_count_47_io_out ? io_r_148_b : _GEN_19127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19129 = 9'h95 == r_count_47_io_out ? io_r_149_b : _GEN_19128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19130 = 9'h96 == r_count_47_io_out ? io_r_150_b : _GEN_19129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19131 = 9'h97 == r_count_47_io_out ? io_r_151_b : _GEN_19130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19132 = 9'h98 == r_count_47_io_out ? io_r_152_b : _GEN_19131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19133 = 9'h99 == r_count_47_io_out ? io_r_153_b : _GEN_19132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19134 = 9'h9a == r_count_47_io_out ? io_r_154_b : _GEN_19133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19135 = 9'h9b == r_count_47_io_out ? io_r_155_b : _GEN_19134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19136 = 9'h9c == r_count_47_io_out ? io_r_156_b : _GEN_19135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19137 = 9'h9d == r_count_47_io_out ? io_r_157_b : _GEN_19136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19138 = 9'h9e == r_count_47_io_out ? io_r_158_b : _GEN_19137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19139 = 9'h9f == r_count_47_io_out ? io_r_159_b : _GEN_19138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19140 = 9'ha0 == r_count_47_io_out ? io_r_160_b : _GEN_19139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19141 = 9'ha1 == r_count_47_io_out ? io_r_161_b : _GEN_19140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19142 = 9'ha2 == r_count_47_io_out ? io_r_162_b : _GEN_19141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19143 = 9'ha3 == r_count_47_io_out ? io_r_163_b : _GEN_19142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19144 = 9'ha4 == r_count_47_io_out ? io_r_164_b : _GEN_19143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19145 = 9'ha5 == r_count_47_io_out ? io_r_165_b : _GEN_19144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19146 = 9'ha6 == r_count_47_io_out ? io_r_166_b : _GEN_19145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19147 = 9'ha7 == r_count_47_io_out ? io_r_167_b : _GEN_19146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19148 = 9'ha8 == r_count_47_io_out ? io_r_168_b : _GEN_19147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19149 = 9'ha9 == r_count_47_io_out ? io_r_169_b : _GEN_19148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19150 = 9'haa == r_count_47_io_out ? io_r_170_b : _GEN_19149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19151 = 9'hab == r_count_47_io_out ? io_r_171_b : _GEN_19150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19152 = 9'hac == r_count_47_io_out ? io_r_172_b : _GEN_19151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19153 = 9'had == r_count_47_io_out ? io_r_173_b : _GEN_19152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19154 = 9'hae == r_count_47_io_out ? io_r_174_b : _GEN_19153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19155 = 9'haf == r_count_47_io_out ? io_r_175_b : _GEN_19154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19156 = 9'hb0 == r_count_47_io_out ? io_r_176_b : _GEN_19155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19157 = 9'hb1 == r_count_47_io_out ? io_r_177_b : _GEN_19156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19158 = 9'hb2 == r_count_47_io_out ? io_r_178_b : _GEN_19157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19159 = 9'hb3 == r_count_47_io_out ? io_r_179_b : _GEN_19158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19160 = 9'hb4 == r_count_47_io_out ? io_r_180_b : _GEN_19159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19161 = 9'hb5 == r_count_47_io_out ? io_r_181_b : _GEN_19160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19162 = 9'hb6 == r_count_47_io_out ? io_r_182_b : _GEN_19161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19163 = 9'hb7 == r_count_47_io_out ? io_r_183_b : _GEN_19162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19164 = 9'hb8 == r_count_47_io_out ? io_r_184_b : _GEN_19163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19165 = 9'hb9 == r_count_47_io_out ? io_r_185_b : _GEN_19164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19166 = 9'hba == r_count_47_io_out ? io_r_186_b : _GEN_19165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19167 = 9'hbb == r_count_47_io_out ? io_r_187_b : _GEN_19166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19168 = 9'hbc == r_count_47_io_out ? io_r_188_b : _GEN_19167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19169 = 9'hbd == r_count_47_io_out ? io_r_189_b : _GEN_19168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19170 = 9'hbe == r_count_47_io_out ? io_r_190_b : _GEN_19169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19171 = 9'hbf == r_count_47_io_out ? io_r_191_b : _GEN_19170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19172 = 9'hc0 == r_count_47_io_out ? io_r_192_b : _GEN_19171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19173 = 9'hc1 == r_count_47_io_out ? io_r_193_b : _GEN_19172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19174 = 9'hc2 == r_count_47_io_out ? io_r_194_b : _GEN_19173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19175 = 9'hc3 == r_count_47_io_out ? io_r_195_b : _GEN_19174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19176 = 9'hc4 == r_count_47_io_out ? io_r_196_b : _GEN_19175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19177 = 9'hc5 == r_count_47_io_out ? io_r_197_b : _GEN_19176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19178 = 9'hc6 == r_count_47_io_out ? io_r_198_b : _GEN_19177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19179 = 9'hc7 == r_count_47_io_out ? io_r_199_b : _GEN_19178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19180 = 9'hc8 == r_count_47_io_out ? io_r_200_b : _GEN_19179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19181 = 9'hc9 == r_count_47_io_out ? io_r_201_b : _GEN_19180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19182 = 9'hca == r_count_47_io_out ? io_r_202_b : _GEN_19181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19183 = 9'hcb == r_count_47_io_out ? io_r_203_b : _GEN_19182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19184 = 9'hcc == r_count_47_io_out ? io_r_204_b : _GEN_19183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19185 = 9'hcd == r_count_47_io_out ? io_r_205_b : _GEN_19184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19186 = 9'hce == r_count_47_io_out ? io_r_206_b : _GEN_19185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19187 = 9'hcf == r_count_47_io_out ? io_r_207_b : _GEN_19186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19188 = 9'hd0 == r_count_47_io_out ? io_r_208_b : _GEN_19187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19189 = 9'hd1 == r_count_47_io_out ? io_r_209_b : _GEN_19188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19190 = 9'hd2 == r_count_47_io_out ? io_r_210_b : _GEN_19189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19191 = 9'hd3 == r_count_47_io_out ? io_r_211_b : _GEN_19190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19192 = 9'hd4 == r_count_47_io_out ? io_r_212_b : _GEN_19191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19193 = 9'hd5 == r_count_47_io_out ? io_r_213_b : _GEN_19192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19194 = 9'hd6 == r_count_47_io_out ? io_r_214_b : _GEN_19193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19195 = 9'hd7 == r_count_47_io_out ? io_r_215_b : _GEN_19194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19196 = 9'hd8 == r_count_47_io_out ? io_r_216_b : _GEN_19195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19197 = 9'hd9 == r_count_47_io_out ? io_r_217_b : _GEN_19196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19198 = 9'hda == r_count_47_io_out ? io_r_218_b : _GEN_19197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19199 = 9'hdb == r_count_47_io_out ? io_r_219_b : _GEN_19198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19200 = 9'hdc == r_count_47_io_out ? io_r_220_b : _GEN_19199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19201 = 9'hdd == r_count_47_io_out ? io_r_221_b : _GEN_19200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19202 = 9'hde == r_count_47_io_out ? io_r_222_b : _GEN_19201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19203 = 9'hdf == r_count_47_io_out ? io_r_223_b : _GEN_19202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19204 = 9'he0 == r_count_47_io_out ? io_r_224_b : _GEN_19203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19205 = 9'he1 == r_count_47_io_out ? io_r_225_b : _GEN_19204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19206 = 9'he2 == r_count_47_io_out ? io_r_226_b : _GEN_19205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19207 = 9'he3 == r_count_47_io_out ? io_r_227_b : _GEN_19206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19208 = 9'he4 == r_count_47_io_out ? io_r_228_b : _GEN_19207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19209 = 9'he5 == r_count_47_io_out ? io_r_229_b : _GEN_19208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19210 = 9'he6 == r_count_47_io_out ? io_r_230_b : _GEN_19209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19211 = 9'he7 == r_count_47_io_out ? io_r_231_b : _GEN_19210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19212 = 9'he8 == r_count_47_io_out ? io_r_232_b : _GEN_19211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19213 = 9'he9 == r_count_47_io_out ? io_r_233_b : _GEN_19212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19214 = 9'hea == r_count_47_io_out ? io_r_234_b : _GEN_19213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19215 = 9'heb == r_count_47_io_out ? io_r_235_b : _GEN_19214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19216 = 9'hec == r_count_47_io_out ? io_r_236_b : _GEN_19215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19217 = 9'hed == r_count_47_io_out ? io_r_237_b : _GEN_19216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19218 = 9'hee == r_count_47_io_out ? io_r_238_b : _GEN_19217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19219 = 9'hef == r_count_47_io_out ? io_r_239_b : _GEN_19218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19220 = 9'hf0 == r_count_47_io_out ? io_r_240_b : _GEN_19219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19221 = 9'hf1 == r_count_47_io_out ? io_r_241_b : _GEN_19220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19222 = 9'hf2 == r_count_47_io_out ? io_r_242_b : _GEN_19221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19223 = 9'hf3 == r_count_47_io_out ? io_r_243_b : _GEN_19222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19224 = 9'hf4 == r_count_47_io_out ? io_r_244_b : _GEN_19223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19225 = 9'hf5 == r_count_47_io_out ? io_r_245_b : _GEN_19224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19226 = 9'hf6 == r_count_47_io_out ? io_r_246_b : _GEN_19225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19227 = 9'hf7 == r_count_47_io_out ? io_r_247_b : _GEN_19226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19228 = 9'hf8 == r_count_47_io_out ? io_r_248_b : _GEN_19227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19229 = 9'hf9 == r_count_47_io_out ? io_r_249_b : _GEN_19228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19230 = 9'hfa == r_count_47_io_out ? io_r_250_b : _GEN_19229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19231 = 9'hfb == r_count_47_io_out ? io_r_251_b : _GEN_19230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19232 = 9'hfc == r_count_47_io_out ? io_r_252_b : _GEN_19231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19233 = 9'hfd == r_count_47_io_out ? io_r_253_b : _GEN_19232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19234 = 9'hfe == r_count_47_io_out ? io_r_254_b : _GEN_19233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19235 = 9'hff == r_count_47_io_out ? io_r_255_b : _GEN_19234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19236 = 9'h100 == r_count_47_io_out ? io_r_256_b : _GEN_19235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19237 = 9'h101 == r_count_47_io_out ? io_r_257_b : _GEN_19236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19238 = 9'h102 == r_count_47_io_out ? io_r_258_b : _GEN_19237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19239 = 9'h103 == r_count_47_io_out ? io_r_259_b : _GEN_19238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19240 = 9'h104 == r_count_47_io_out ? io_r_260_b : _GEN_19239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19241 = 9'h105 == r_count_47_io_out ? io_r_261_b : _GEN_19240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19242 = 9'h106 == r_count_47_io_out ? io_r_262_b : _GEN_19241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19243 = 9'h107 == r_count_47_io_out ? io_r_263_b : _GEN_19242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19244 = 9'h108 == r_count_47_io_out ? io_r_264_b : _GEN_19243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19245 = 9'h109 == r_count_47_io_out ? io_r_265_b : _GEN_19244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19246 = 9'h10a == r_count_47_io_out ? io_r_266_b : _GEN_19245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19247 = 9'h10b == r_count_47_io_out ? io_r_267_b : _GEN_19246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19248 = 9'h10c == r_count_47_io_out ? io_r_268_b : _GEN_19247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19249 = 9'h10d == r_count_47_io_out ? io_r_269_b : _GEN_19248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19250 = 9'h10e == r_count_47_io_out ? io_r_270_b : _GEN_19249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19251 = 9'h10f == r_count_47_io_out ? io_r_271_b : _GEN_19250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19252 = 9'h110 == r_count_47_io_out ? io_r_272_b : _GEN_19251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19253 = 9'h111 == r_count_47_io_out ? io_r_273_b : _GEN_19252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19254 = 9'h112 == r_count_47_io_out ? io_r_274_b : _GEN_19253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19255 = 9'h113 == r_count_47_io_out ? io_r_275_b : _GEN_19254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19256 = 9'h114 == r_count_47_io_out ? io_r_276_b : _GEN_19255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19257 = 9'h115 == r_count_47_io_out ? io_r_277_b : _GEN_19256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19258 = 9'h116 == r_count_47_io_out ? io_r_278_b : _GEN_19257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19259 = 9'h117 == r_count_47_io_out ? io_r_279_b : _GEN_19258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19260 = 9'h118 == r_count_47_io_out ? io_r_280_b : _GEN_19259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19261 = 9'h119 == r_count_47_io_out ? io_r_281_b : _GEN_19260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19262 = 9'h11a == r_count_47_io_out ? io_r_282_b : _GEN_19261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19263 = 9'h11b == r_count_47_io_out ? io_r_283_b : _GEN_19262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19264 = 9'h11c == r_count_47_io_out ? io_r_284_b : _GEN_19263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19265 = 9'h11d == r_count_47_io_out ? io_r_285_b : _GEN_19264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19266 = 9'h11e == r_count_47_io_out ? io_r_286_b : _GEN_19265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19267 = 9'h11f == r_count_47_io_out ? io_r_287_b : _GEN_19266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19268 = 9'h120 == r_count_47_io_out ? io_r_288_b : _GEN_19267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19269 = 9'h121 == r_count_47_io_out ? io_r_289_b : _GEN_19268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19270 = 9'h122 == r_count_47_io_out ? io_r_290_b : _GEN_19269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19271 = 9'h123 == r_count_47_io_out ? io_r_291_b : _GEN_19270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19272 = 9'h124 == r_count_47_io_out ? io_r_292_b : _GEN_19271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19273 = 9'h125 == r_count_47_io_out ? io_r_293_b : _GEN_19272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19274 = 9'h126 == r_count_47_io_out ? io_r_294_b : _GEN_19273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19275 = 9'h127 == r_count_47_io_out ? io_r_295_b : _GEN_19274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19276 = 9'h128 == r_count_47_io_out ? io_r_296_b : _GEN_19275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19277 = 9'h129 == r_count_47_io_out ? io_r_297_b : _GEN_19276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19278 = 9'h12a == r_count_47_io_out ? io_r_298_b : _GEN_19277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19279 = 9'h12b == r_count_47_io_out ? io_r_299_b : _GEN_19278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19280 = 9'h12c == r_count_47_io_out ? io_r_300_b : _GEN_19279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19281 = 9'h12d == r_count_47_io_out ? io_r_301_b : _GEN_19280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19282 = 9'h12e == r_count_47_io_out ? io_r_302_b : _GEN_19281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19283 = 9'h12f == r_count_47_io_out ? io_r_303_b : _GEN_19282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19284 = 9'h130 == r_count_47_io_out ? io_r_304_b : _GEN_19283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19285 = 9'h131 == r_count_47_io_out ? io_r_305_b : _GEN_19284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19286 = 9'h132 == r_count_47_io_out ? io_r_306_b : _GEN_19285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19287 = 9'h133 == r_count_47_io_out ? io_r_307_b : _GEN_19286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19288 = 9'h134 == r_count_47_io_out ? io_r_308_b : _GEN_19287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19289 = 9'h135 == r_count_47_io_out ? io_r_309_b : _GEN_19288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19290 = 9'h136 == r_count_47_io_out ? io_r_310_b : _GEN_19289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19291 = 9'h137 == r_count_47_io_out ? io_r_311_b : _GEN_19290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19292 = 9'h138 == r_count_47_io_out ? io_r_312_b : _GEN_19291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19293 = 9'h139 == r_count_47_io_out ? io_r_313_b : _GEN_19292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19294 = 9'h13a == r_count_47_io_out ? io_r_314_b : _GEN_19293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19295 = 9'h13b == r_count_47_io_out ? io_r_315_b : _GEN_19294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19296 = 9'h13c == r_count_47_io_out ? io_r_316_b : _GEN_19295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19297 = 9'h13d == r_count_47_io_out ? io_r_317_b : _GEN_19296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19298 = 9'h13e == r_count_47_io_out ? io_r_318_b : _GEN_19297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19299 = 9'h13f == r_count_47_io_out ? io_r_319_b : _GEN_19298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19300 = 9'h140 == r_count_47_io_out ? io_r_320_b : _GEN_19299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19301 = 9'h141 == r_count_47_io_out ? io_r_321_b : _GEN_19300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19302 = 9'h142 == r_count_47_io_out ? io_r_322_b : _GEN_19301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19303 = 9'h143 == r_count_47_io_out ? io_r_323_b : _GEN_19302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19304 = 9'h144 == r_count_47_io_out ? io_r_324_b : _GEN_19303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19305 = 9'h145 == r_count_47_io_out ? io_r_325_b : _GEN_19304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19306 = 9'h146 == r_count_47_io_out ? io_r_326_b : _GEN_19305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19307 = 9'h147 == r_count_47_io_out ? io_r_327_b : _GEN_19306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19308 = 9'h148 == r_count_47_io_out ? io_r_328_b : _GEN_19307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19309 = 9'h149 == r_count_47_io_out ? io_r_329_b : _GEN_19308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19310 = 9'h14a == r_count_47_io_out ? io_r_330_b : _GEN_19309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19311 = 9'h14b == r_count_47_io_out ? io_r_331_b : _GEN_19310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19312 = 9'h14c == r_count_47_io_out ? io_r_332_b : _GEN_19311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19313 = 9'h14d == r_count_47_io_out ? io_r_333_b : _GEN_19312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19314 = 9'h14e == r_count_47_io_out ? io_r_334_b : _GEN_19313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19315 = 9'h14f == r_count_47_io_out ? io_r_335_b : _GEN_19314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19316 = 9'h150 == r_count_47_io_out ? io_r_336_b : _GEN_19315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19317 = 9'h151 == r_count_47_io_out ? io_r_337_b : _GEN_19316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19318 = 9'h152 == r_count_47_io_out ? io_r_338_b : _GEN_19317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19319 = 9'h153 == r_count_47_io_out ? io_r_339_b : _GEN_19318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19320 = 9'h154 == r_count_47_io_out ? io_r_340_b : _GEN_19319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19321 = 9'h155 == r_count_47_io_out ? io_r_341_b : _GEN_19320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19322 = 9'h156 == r_count_47_io_out ? io_r_342_b : _GEN_19321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19323 = 9'h157 == r_count_47_io_out ? io_r_343_b : _GEN_19322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19324 = 9'h158 == r_count_47_io_out ? io_r_344_b : _GEN_19323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19325 = 9'h159 == r_count_47_io_out ? io_r_345_b : _GEN_19324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19326 = 9'h15a == r_count_47_io_out ? io_r_346_b : _GEN_19325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19327 = 9'h15b == r_count_47_io_out ? io_r_347_b : _GEN_19326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19328 = 9'h15c == r_count_47_io_out ? io_r_348_b : _GEN_19327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19329 = 9'h15d == r_count_47_io_out ? io_r_349_b : _GEN_19328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19330 = 9'h15e == r_count_47_io_out ? io_r_350_b : _GEN_19329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19331 = 9'h15f == r_count_47_io_out ? io_r_351_b : _GEN_19330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19332 = 9'h160 == r_count_47_io_out ? io_r_352_b : _GEN_19331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19333 = 9'h161 == r_count_47_io_out ? io_r_353_b : _GEN_19332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19334 = 9'h162 == r_count_47_io_out ? io_r_354_b : _GEN_19333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19335 = 9'h163 == r_count_47_io_out ? io_r_355_b : _GEN_19334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19336 = 9'h164 == r_count_47_io_out ? io_r_356_b : _GEN_19335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19337 = 9'h165 == r_count_47_io_out ? io_r_357_b : _GEN_19336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19338 = 9'h166 == r_count_47_io_out ? io_r_358_b : _GEN_19337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19339 = 9'h167 == r_count_47_io_out ? io_r_359_b : _GEN_19338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19340 = 9'h168 == r_count_47_io_out ? io_r_360_b : _GEN_19339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19341 = 9'h169 == r_count_47_io_out ? io_r_361_b : _GEN_19340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19342 = 9'h16a == r_count_47_io_out ? io_r_362_b : _GEN_19341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19343 = 9'h16b == r_count_47_io_out ? io_r_363_b : _GEN_19342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19344 = 9'h16c == r_count_47_io_out ? io_r_364_b : _GEN_19343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19345 = 9'h16d == r_count_47_io_out ? io_r_365_b : _GEN_19344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19346 = 9'h16e == r_count_47_io_out ? io_r_366_b : _GEN_19345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19347 = 9'h16f == r_count_47_io_out ? io_r_367_b : _GEN_19346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19348 = 9'h170 == r_count_47_io_out ? io_r_368_b : _GEN_19347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19349 = 9'h171 == r_count_47_io_out ? io_r_369_b : _GEN_19348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19350 = 9'h172 == r_count_47_io_out ? io_r_370_b : _GEN_19349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19351 = 9'h173 == r_count_47_io_out ? io_r_371_b : _GEN_19350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19352 = 9'h174 == r_count_47_io_out ? io_r_372_b : _GEN_19351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19353 = 9'h175 == r_count_47_io_out ? io_r_373_b : _GEN_19352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19354 = 9'h176 == r_count_47_io_out ? io_r_374_b : _GEN_19353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19355 = 9'h177 == r_count_47_io_out ? io_r_375_b : _GEN_19354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19356 = 9'h178 == r_count_47_io_out ? io_r_376_b : _GEN_19355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19357 = 9'h179 == r_count_47_io_out ? io_r_377_b : _GEN_19356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19358 = 9'h17a == r_count_47_io_out ? io_r_378_b : _GEN_19357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19359 = 9'h17b == r_count_47_io_out ? io_r_379_b : _GEN_19358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19360 = 9'h17c == r_count_47_io_out ? io_r_380_b : _GEN_19359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19361 = 9'h17d == r_count_47_io_out ? io_r_381_b : _GEN_19360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19362 = 9'h17e == r_count_47_io_out ? io_r_382_b : _GEN_19361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19363 = 9'h17f == r_count_47_io_out ? io_r_383_b : _GEN_19362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19364 = 9'h180 == r_count_47_io_out ? io_r_384_b : _GEN_19363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19365 = 9'h181 == r_count_47_io_out ? io_r_385_b : _GEN_19364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19366 = 9'h182 == r_count_47_io_out ? io_r_386_b : _GEN_19365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19367 = 9'h183 == r_count_47_io_out ? io_r_387_b : _GEN_19366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19368 = 9'h184 == r_count_47_io_out ? io_r_388_b : _GEN_19367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19369 = 9'h185 == r_count_47_io_out ? io_r_389_b : _GEN_19368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19370 = 9'h186 == r_count_47_io_out ? io_r_390_b : _GEN_19369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19371 = 9'h187 == r_count_47_io_out ? io_r_391_b : _GEN_19370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19372 = 9'h188 == r_count_47_io_out ? io_r_392_b : _GEN_19371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19373 = 9'h189 == r_count_47_io_out ? io_r_393_b : _GEN_19372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19374 = 9'h18a == r_count_47_io_out ? io_r_394_b : _GEN_19373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19375 = 9'h18b == r_count_47_io_out ? io_r_395_b : _GEN_19374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19376 = 9'h18c == r_count_47_io_out ? io_r_396_b : _GEN_19375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19377 = 9'h18d == r_count_47_io_out ? io_r_397_b : _GEN_19376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19378 = 9'h18e == r_count_47_io_out ? io_r_398_b : _GEN_19377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19381 = 9'h1 == r_count_48_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19382 = 9'h2 == r_count_48_io_out ? io_r_2_b : _GEN_19381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19383 = 9'h3 == r_count_48_io_out ? io_r_3_b : _GEN_19382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19384 = 9'h4 == r_count_48_io_out ? io_r_4_b : _GEN_19383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19385 = 9'h5 == r_count_48_io_out ? io_r_5_b : _GEN_19384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19386 = 9'h6 == r_count_48_io_out ? io_r_6_b : _GEN_19385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19387 = 9'h7 == r_count_48_io_out ? io_r_7_b : _GEN_19386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19388 = 9'h8 == r_count_48_io_out ? io_r_8_b : _GEN_19387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19389 = 9'h9 == r_count_48_io_out ? io_r_9_b : _GEN_19388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19390 = 9'ha == r_count_48_io_out ? io_r_10_b : _GEN_19389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19391 = 9'hb == r_count_48_io_out ? io_r_11_b : _GEN_19390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19392 = 9'hc == r_count_48_io_out ? io_r_12_b : _GEN_19391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19393 = 9'hd == r_count_48_io_out ? io_r_13_b : _GEN_19392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19394 = 9'he == r_count_48_io_out ? io_r_14_b : _GEN_19393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19395 = 9'hf == r_count_48_io_out ? io_r_15_b : _GEN_19394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19396 = 9'h10 == r_count_48_io_out ? io_r_16_b : _GEN_19395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19397 = 9'h11 == r_count_48_io_out ? io_r_17_b : _GEN_19396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19398 = 9'h12 == r_count_48_io_out ? io_r_18_b : _GEN_19397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19399 = 9'h13 == r_count_48_io_out ? io_r_19_b : _GEN_19398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19400 = 9'h14 == r_count_48_io_out ? io_r_20_b : _GEN_19399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19401 = 9'h15 == r_count_48_io_out ? io_r_21_b : _GEN_19400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19402 = 9'h16 == r_count_48_io_out ? io_r_22_b : _GEN_19401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19403 = 9'h17 == r_count_48_io_out ? io_r_23_b : _GEN_19402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19404 = 9'h18 == r_count_48_io_out ? io_r_24_b : _GEN_19403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19405 = 9'h19 == r_count_48_io_out ? io_r_25_b : _GEN_19404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19406 = 9'h1a == r_count_48_io_out ? io_r_26_b : _GEN_19405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19407 = 9'h1b == r_count_48_io_out ? io_r_27_b : _GEN_19406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19408 = 9'h1c == r_count_48_io_out ? io_r_28_b : _GEN_19407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19409 = 9'h1d == r_count_48_io_out ? io_r_29_b : _GEN_19408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19410 = 9'h1e == r_count_48_io_out ? io_r_30_b : _GEN_19409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19411 = 9'h1f == r_count_48_io_out ? io_r_31_b : _GEN_19410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19412 = 9'h20 == r_count_48_io_out ? io_r_32_b : _GEN_19411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19413 = 9'h21 == r_count_48_io_out ? io_r_33_b : _GEN_19412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19414 = 9'h22 == r_count_48_io_out ? io_r_34_b : _GEN_19413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19415 = 9'h23 == r_count_48_io_out ? io_r_35_b : _GEN_19414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19416 = 9'h24 == r_count_48_io_out ? io_r_36_b : _GEN_19415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19417 = 9'h25 == r_count_48_io_out ? io_r_37_b : _GEN_19416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19418 = 9'h26 == r_count_48_io_out ? io_r_38_b : _GEN_19417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19419 = 9'h27 == r_count_48_io_out ? io_r_39_b : _GEN_19418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19420 = 9'h28 == r_count_48_io_out ? io_r_40_b : _GEN_19419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19421 = 9'h29 == r_count_48_io_out ? io_r_41_b : _GEN_19420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19422 = 9'h2a == r_count_48_io_out ? io_r_42_b : _GEN_19421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19423 = 9'h2b == r_count_48_io_out ? io_r_43_b : _GEN_19422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19424 = 9'h2c == r_count_48_io_out ? io_r_44_b : _GEN_19423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19425 = 9'h2d == r_count_48_io_out ? io_r_45_b : _GEN_19424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19426 = 9'h2e == r_count_48_io_out ? io_r_46_b : _GEN_19425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19427 = 9'h2f == r_count_48_io_out ? io_r_47_b : _GEN_19426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19428 = 9'h30 == r_count_48_io_out ? io_r_48_b : _GEN_19427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19429 = 9'h31 == r_count_48_io_out ? io_r_49_b : _GEN_19428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19430 = 9'h32 == r_count_48_io_out ? io_r_50_b : _GEN_19429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19431 = 9'h33 == r_count_48_io_out ? io_r_51_b : _GEN_19430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19432 = 9'h34 == r_count_48_io_out ? io_r_52_b : _GEN_19431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19433 = 9'h35 == r_count_48_io_out ? io_r_53_b : _GEN_19432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19434 = 9'h36 == r_count_48_io_out ? io_r_54_b : _GEN_19433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19435 = 9'h37 == r_count_48_io_out ? io_r_55_b : _GEN_19434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19436 = 9'h38 == r_count_48_io_out ? io_r_56_b : _GEN_19435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19437 = 9'h39 == r_count_48_io_out ? io_r_57_b : _GEN_19436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19438 = 9'h3a == r_count_48_io_out ? io_r_58_b : _GEN_19437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19439 = 9'h3b == r_count_48_io_out ? io_r_59_b : _GEN_19438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19440 = 9'h3c == r_count_48_io_out ? io_r_60_b : _GEN_19439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19441 = 9'h3d == r_count_48_io_out ? io_r_61_b : _GEN_19440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19442 = 9'h3e == r_count_48_io_out ? io_r_62_b : _GEN_19441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19443 = 9'h3f == r_count_48_io_out ? io_r_63_b : _GEN_19442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19444 = 9'h40 == r_count_48_io_out ? io_r_64_b : _GEN_19443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19445 = 9'h41 == r_count_48_io_out ? io_r_65_b : _GEN_19444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19446 = 9'h42 == r_count_48_io_out ? io_r_66_b : _GEN_19445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19447 = 9'h43 == r_count_48_io_out ? io_r_67_b : _GEN_19446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19448 = 9'h44 == r_count_48_io_out ? io_r_68_b : _GEN_19447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19449 = 9'h45 == r_count_48_io_out ? io_r_69_b : _GEN_19448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19450 = 9'h46 == r_count_48_io_out ? io_r_70_b : _GEN_19449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19451 = 9'h47 == r_count_48_io_out ? io_r_71_b : _GEN_19450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19452 = 9'h48 == r_count_48_io_out ? io_r_72_b : _GEN_19451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19453 = 9'h49 == r_count_48_io_out ? io_r_73_b : _GEN_19452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19454 = 9'h4a == r_count_48_io_out ? io_r_74_b : _GEN_19453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19455 = 9'h4b == r_count_48_io_out ? io_r_75_b : _GEN_19454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19456 = 9'h4c == r_count_48_io_out ? io_r_76_b : _GEN_19455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19457 = 9'h4d == r_count_48_io_out ? io_r_77_b : _GEN_19456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19458 = 9'h4e == r_count_48_io_out ? io_r_78_b : _GEN_19457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19459 = 9'h4f == r_count_48_io_out ? io_r_79_b : _GEN_19458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19460 = 9'h50 == r_count_48_io_out ? io_r_80_b : _GEN_19459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19461 = 9'h51 == r_count_48_io_out ? io_r_81_b : _GEN_19460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19462 = 9'h52 == r_count_48_io_out ? io_r_82_b : _GEN_19461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19463 = 9'h53 == r_count_48_io_out ? io_r_83_b : _GEN_19462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19464 = 9'h54 == r_count_48_io_out ? io_r_84_b : _GEN_19463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19465 = 9'h55 == r_count_48_io_out ? io_r_85_b : _GEN_19464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19466 = 9'h56 == r_count_48_io_out ? io_r_86_b : _GEN_19465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19467 = 9'h57 == r_count_48_io_out ? io_r_87_b : _GEN_19466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19468 = 9'h58 == r_count_48_io_out ? io_r_88_b : _GEN_19467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19469 = 9'h59 == r_count_48_io_out ? io_r_89_b : _GEN_19468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19470 = 9'h5a == r_count_48_io_out ? io_r_90_b : _GEN_19469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19471 = 9'h5b == r_count_48_io_out ? io_r_91_b : _GEN_19470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19472 = 9'h5c == r_count_48_io_out ? io_r_92_b : _GEN_19471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19473 = 9'h5d == r_count_48_io_out ? io_r_93_b : _GEN_19472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19474 = 9'h5e == r_count_48_io_out ? io_r_94_b : _GEN_19473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19475 = 9'h5f == r_count_48_io_out ? io_r_95_b : _GEN_19474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19476 = 9'h60 == r_count_48_io_out ? io_r_96_b : _GEN_19475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19477 = 9'h61 == r_count_48_io_out ? io_r_97_b : _GEN_19476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19478 = 9'h62 == r_count_48_io_out ? io_r_98_b : _GEN_19477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19479 = 9'h63 == r_count_48_io_out ? io_r_99_b : _GEN_19478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19480 = 9'h64 == r_count_48_io_out ? io_r_100_b : _GEN_19479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19481 = 9'h65 == r_count_48_io_out ? io_r_101_b : _GEN_19480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19482 = 9'h66 == r_count_48_io_out ? io_r_102_b : _GEN_19481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19483 = 9'h67 == r_count_48_io_out ? io_r_103_b : _GEN_19482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19484 = 9'h68 == r_count_48_io_out ? io_r_104_b : _GEN_19483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19485 = 9'h69 == r_count_48_io_out ? io_r_105_b : _GEN_19484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19486 = 9'h6a == r_count_48_io_out ? io_r_106_b : _GEN_19485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19487 = 9'h6b == r_count_48_io_out ? io_r_107_b : _GEN_19486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19488 = 9'h6c == r_count_48_io_out ? io_r_108_b : _GEN_19487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19489 = 9'h6d == r_count_48_io_out ? io_r_109_b : _GEN_19488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19490 = 9'h6e == r_count_48_io_out ? io_r_110_b : _GEN_19489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19491 = 9'h6f == r_count_48_io_out ? io_r_111_b : _GEN_19490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19492 = 9'h70 == r_count_48_io_out ? io_r_112_b : _GEN_19491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19493 = 9'h71 == r_count_48_io_out ? io_r_113_b : _GEN_19492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19494 = 9'h72 == r_count_48_io_out ? io_r_114_b : _GEN_19493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19495 = 9'h73 == r_count_48_io_out ? io_r_115_b : _GEN_19494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19496 = 9'h74 == r_count_48_io_out ? io_r_116_b : _GEN_19495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19497 = 9'h75 == r_count_48_io_out ? io_r_117_b : _GEN_19496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19498 = 9'h76 == r_count_48_io_out ? io_r_118_b : _GEN_19497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19499 = 9'h77 == r_count_48_io_out ? io_r_119_b : _GEN_19498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19500 = 9'h78 == r_count_48_io_out ? io_r_120_b : _GEN_19499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19501 = 9'h79 == r_count_48_io_out ? io_r_121_b : _GEN_19500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19502 = 9'h7a == r_count_48_io_out ? io_r_122_b : _GEN_19501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19503 = 9'h7b == r_count_48_io_out ? io_r_123_b : _GEN_19502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19504 = 9'h7c == r_count_48_io_out ? io_r_124_b : _GEN_19503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19505 = 9'h7d == r_count_48_io_out ? io_r_125_b : _GEN_19504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19506 = 9'h7e == r_count_48_io_out ? io_r_126_b : _GEN_19505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19507 = 9'h7f == r_count_48_io_out ? io_r_127_b : _GEN_19506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19508 = 9'h80 == r_count_48_io_out ? io_r_128_b : _GEN_19507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19509 = 9'h81 == r_count_48_io_out ? io_r_129_b : _GEN_19508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19510 = 9'h82 == r_count_48_io_out ? io_r_130_b : _GEN_19509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19511 = 9'h83 == r_count_48_io_out ? io_r_131_b : _GEN_19510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19512 = 9'h84 == r_count_48_io_out ? io_r_132_b : _GEN_19511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19513 = 9'h85 == r_count_48_io_out ? io_r_133_b : _GEN_19512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19514 = 9'h86 == r_count_48_io_out ? io_r_134_b : _GEN_19513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19515 = 9'h87 == r_count_48_io_out ? io_r_135_b : _GEN_19514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19516 = 9'h88 == r_count_48_io_out ? io_r_136_b : _GEN_19515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19517 = 9'h89 == r_count_48_io_out ? io_r_137_b : _GEN_19516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19518 = 9'h8a == r_count_48_io_out ? io_r_138_b : _GEN_19517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19519 = 9'h8b == r_count_48_io_out ? io_r_139_b : _GEN_19518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19520 = 9'h8c == r_count_48_io_out ? io_r_140_b : _GEN_19519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19521 = 9'h8d == r_count_48_io_out ? io_r_141_b : _GEN_19520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19522 = 9'h8e == r_count_48_io_out ? io_r_142_b : _GEN_19521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19523 = 9'h8f == r_count_48_io_out ? io_r_143_b : _GEN_19522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19524 = 9'h90 == r_count_48_io_out ? io_r_144_b : _GEN_19523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19525 = 9'h91 == r_count_48_io_out ? io_r_145_b : _GEN_19524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19526 = 9'h92 == r_count_48_io_out ? io_r_146_b : _GEN_19525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19527 = 9'h93 == r_count_48_io_out ? io_r_147_b : _GEN_19526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19528 = 9'h94 == r_count_48_io_out ? io_r_148_b : _GEN_19527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19529 = 9'h95 == r_count_48_io_out ? io_r_149_b : _GEN_19528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19530 = 9'h96 == r_count_48_io_out ? io_r_150_b : _GEN_19529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19531 = 9'h97 == r_count_48_io_out ? io_r_151_b : _GEN_19530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19532 = 9'h98 == r_count_48_io_out ? io_r_152_b : _GEN_19531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19533 = 9'h99 == r_count_48_io_out ? io_r_153_b : _GEN_19532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19534 = 9'h9a == r_count_48_io_out ? io_r_154_b : _GEN_19533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19535 = 9'h9b == r_count_48_io_out ? io_r_155_b : _GEN_19534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19536 = 9'h9c == r_count_48_io_out ? io_r_156_b : _GEN_19535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19537 = 9'h9d == r_count_48_io_out ? io_r_157_b : _GEN_19536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19538 = 9'h9e == r_count_48_io_out ? io_r_158_b : _GEN_19537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19539 = 9'h9f == r_count_48_io_out ? io_r_159_b : _GEN_19538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19540 = 9'ha0 == r_count_48_io_out ? io_r_160_b : _GEN_19539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19541 = 9'ha1 == r_count_48_io_out ? io_r_161_b : _GEN_19540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19542 = 9'ha2 == r_count_48_io_out ? io_r_162_b : _GEN_19541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19543 = 9'ha3 == r_count_48_io_out ? io_r_163_b : _GEN_19542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19544 = 9'ha4 == r_count_48_io_out ? io_r_164_b : _GEN_19543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19545 = 9'ha5 == r_count_48_io_out ? io_r_165_b : _GEN_19544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19546 = 9'ha6 == r_count_48_io_out ? io_r_166_b : _GEN_19545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19547 = 9'ha7 == r_count_48_io_out ? io_r_167_b : _GEN_19546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19548 = 9'ha8 == r_count_48_io_out ? io_r_168_b : _GEN_19547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19549 = 9'ha9 == r_count_48_io_out ? io_r_169_b : _GEN_19548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19550 = 9'haa == r_count_48_io_out ? io_r_170_b : _GEN_19549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19551 = 9'hab == r_count_48_io_out ? io_r_171_b : _GEN_19550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19552 = 9'hac == r_count_48_io_out ? io_r_172_b : _GEN_19551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19553 = 9'had == r_count_48_io_out ? io_r_173_b : _GEN_19552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19554 = 9'hae == r_count_48_io_out ? io_r_174_b : _GEN_19553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19555 = 9'haf == r_count_48_io_out ? io_r_175_b : _GEN_19554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19556 = 9'hb0 == r_count_48_io_out ? io_r_176_b : _GEN_19555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19557 = 9'hb1 == r_count_48_io_out ? io_r_177_b : _GEN_19556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19558 = 9'hb2 == r_count_48_io_out ? io_r_178_b : _GEN_19557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19559 = 9'hb3 == r_count_48_io_out ? io_r_179_b : _GEN_19558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19560 = 9'hb4 == r_count_48_io_out ? io_r_180_b : _GEN_19559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19561 = 9'hb5 == r_count_48_io_out ? io_r_181_b : _GEN_19560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19562 = 9'hb6 == r_count_48_io_out ? io_r_182_b : _GEN_19561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19563 = 9'hb7 == r_count_48_io_out ? io_r_183_b : _GEN_19562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19564 = 9'hb8 == r_count_48_io_out ? io_r_184_b : _GEN_19563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19565 = 9'hb9 == r_count_48_io_out ? io_r_185_b : _GEN_19564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19566 = 9'hba == r_count_48_io_out ? io_r_186_b : _GEN_19565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19567 = 9'hbb == r_count_48_io_out ? io_r_187_b : _GEN_19566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19568 = 9'hbc == r_count_48_io_out ? io_r_188_b : _GEN_19567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19569 = 9'hbd == r_count_48_io_out ? io_r_189_b : _GEN_19568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19570 = 9'hbe == r_count_48_io_out ? io_r_190_b : _GEN_19569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19571 = 9'hbf == r_count_48_io_out ? io_r_191_b : _GEN_19570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19572 = 9'hc0 == r_count_48_io_out ? io_r_192_b : _GEN_19571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19573 = 9'hc1 == r_count_48_io_out ? io_r_193_b : _GEN_19572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19574 = 9'hc2 == r_count_48_io_out ? io_r_194_b : _GEN_19573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19575 = 9'hc3 == r_count_48_io_out ? io_r_195_b : _GEN_19574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19576 = 9'hc4 == r_count_48_io_out ? io_r_196_b : _GEN_19575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19577 = 9'hc5 == r_count_48_io_out ? io_r_197_b : _GEN_19576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19578 = 9'hc6 == r_count_48_io_out ? io_r_198_b : _GEN_19577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19579 = 9'hc7 == r_count_48_io_out ? io_r_199_b : _GEN_19578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19580 = 9'hc8 == r_count_48_io_out ? io_r_200_b : _GEN_19579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19581 = 9'hc9 == r_count_48_io_out ? io_r_201_b : _GEN_19580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19582 = 9'hca == r_count_48_io_out ? io_r_202_b : _GEN_19581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19583 = 9'hcb == r_count_48_io_out ? io_r_203_b : _GEN_19582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19584 = 9'hcc == r_count_48_io_out ? io_r_204_b : _GEN_19583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19585 = 9'hcd == r_count_48_io_out ? io_r_205_b : _GEN_19584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19586 = 9'hce == r_count_48_io_out ? io_r_206_b : _GEN_19585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19587 = 9'hcf == r_count_48_io_out ? io_r_207_b : _GEN_19586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19588 = 9'hd0 == r_count_48_io_out ? io_r_208_b : _GEN_19587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19589 = 9'hd1 == r_count_48_io_out ? io_r_209_b : _GEN_19588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19590 = 9'hd2 == r_count_48_io_out ? io_r_210_b : _GEN_19589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19591 = 9'hd3 == r_count_48_io_out ? io_r_211_b : _GEN_19590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19592 = 9'hd4 == r_count_48_io_out ? io_r_212_b : _GEN_19591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19593 = 9'hd5 == r_count_48_io_out ? io_r_213_b : _GEN_19592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19594 = 9'hd6 == r_count_48_io_out ? io_r_214_b : _GEN_19593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19595 = 9'hd7 == r_count_48_io_out ? io_r_215_b : _GEN_19594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19596 = 9'hd8 == r_count_48_io_out ? io_r_216_b : _GEN_19595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19597 = 9'hd9 == r_count_48_io_out ? io_r_217_b : _GEN_19596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19598 = 9'hda == r_count_48_io_out ? io_r_218_b : _GEN_19597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19599 = 9'hdb == r_count_48_io_out ? io_r_219_b : _GEN_19598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19600 = 9'hdc == r_count_48_io_out ? io_r_220_b : _GEN_19599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19601 = 9'hdd == r_count_48_io_out ? io_r_221_b : _GEN_19600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19602 = 9'hde == r_count_48_io_out ? io_r_222_b : _GEN_19601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19603 = 9'hdf == r_count_48_io_out ? io_r_223_b : _GEN_19602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19604 = 9'he0 == r_count_48_io_out ? io_r_224_b : _GEN_19603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19605 = 9'he1 == r_count_48_io_out ? io_r_225_b : _GEN_19604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19606 = 9'he2 == r_count_48_io_out ? io_r_226_b : _GEN_19605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19607 = 9'he3 == r_count_48_io_out ? io_r_227_b : _GEN_19606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19608 = 9'he4 == r_count_48_io_out ? io_r_228_b : _GEN_19607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19609 = 9'he5 == r_count_48_io_out ? io_r_229_b : _GEN_19608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19610 = 9'he6 == r_count_48_io_out ? io_r_230_b : _GEN_19609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19611 = 9'he7 == r_count_48_io_out ? io_r_231_b : _GEN_19610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19612 = 9'he8 == r_count_48_io_out ? io_r_232_b : _GEN_19611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19613 = 9'he9 == r_count_48_io_out ? io_r_233_b : _GEN_19612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19614 = 9'hea == r_count_48_io_out ? io_r_234_b : _GEN_19613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19615 = 9'heb == r_count_48_io_out ? io_r_235_b : _GEN_19614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19616 = 9'hec == r_count_48_io_out ? io_r_236_b : _GEN_19615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19617 = 9'hed == r_count_48_io_out ? io_r_237_b : _GEN_19616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19618 = 9'hee == r_count_48_io_out ? io_r_238_b : _GEN_19617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19619 = 9'hef == r_count_48_io_out ? io_r_239_b : _GEN_19618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19620 = 9'hf0 == r_count_48_io_out ? io_r_240_b : _GEN_19619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19621 = 9'hf1 == r_count_48_io_out ? io_r_241_b : _GEN_19620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19622 = 9'hf2 == r_count_48_io_out ? io_r_242_b : _GEN_19621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19623 = 9'hf3 == r_count_48_io_out ? io_r_243_b : _GEN_19622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19624 = 9'hf4 == r_count_48_io_out ? io_r_244_b : _GEN_19623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19625 = 9'hf5 == r_count_48_io_out ? io_r_245_b : _GEN_19624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19626 = 9'hf6 == r_count_48_io_out ? io_r_246_b : _GEN_19625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19627 = 9'hf7 == r_count_48_io_out ? io_r_247_b : _GEN_19626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19628 = 9'hf8 == r_count_48_io_out ? io_r_248_b : _GEN_19627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19629 = 9'hf9 == r_count_48_io_out ? io_r_249_b : _GEN_19628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19630 = 9'hfa == r_count_48_io_out ? io_r_250_b : _GEN_19629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19631 = 9'hfb == r_count_48_io_out ? io_r_251_b : _GEN_19630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19632 = 9'hfc == r_count_48_io_out ? io_r_252_b : _GEN_19631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19633 = 9'hfd == r_count_48_io_out ? io_r_253_b : _GEN_19632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19634 = 9'hfe == r_count_48_io_out ? io_r_254_b : _GEN_19633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19635 = 9'hff == r_count_48_io_out ? io_r_255_b : _GEN_19634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19636 = 9'h100 == r_count_48_io_out ? io_r_256_b : _GEN_19635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19637 = 9'h101 == r_count_48_io_out ? io_r_257_b : _GEN_19636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19638 = 9'h102 == r_count_48_io_out ? io_r_258_b : _GEN_19637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19639 = 9'h103 == r_count_48_io_out ? io_r_259_b : _GEN_19638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19640 = 9'h104 == r_count_48_io_out ? io_r_260_b : _GEN_19639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19641 = 9'h105 == r_count_48_io_out ? io_r_261_b : _GEN_19640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19642 = 9'h106 == r_count_48_io_out ? io_r_262_b : _GEN_19641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19643 = 9'h107 == r_count_48_io_out ? io_r_263_b : _GEN_19642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19644 = 9'h108 == r_count_48_io_out ? io_r_264_b : _GEN_19643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19645 = 9'h109 == r_count_48_io_out ? io_r_265_b : _GEN_19644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19646 = 9'h10a == r_count_48_io_out ? io_r_266_b : _GEN_19645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19647 = 9'h10b == r_count_48_io_out ? io_r_267_b : _GEN_19646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19648 = 9'h10c == r_count_48_io_out ? io_r_268_b : _GEN_19647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19649 = 9'h10d == r_count_48_io_out ? io_r_269_b : _GEN_19648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19650 = 9'h10e == r_count_48_io_out ? io_r_270_b : _GEN_19649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19651 = 9'h10f == r_count_48_io_out ? io_r_271_b : _GEN_19650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19652 = 9'h110 == r_count_48_io_out ? io_r_272_b : _GEN_19651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19653 = 9'h111 == r_count_48_io_out ? io_r_273_b : _GEN_19652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19654 = 9'h112 == r_count_48_io_out ? io_r_274_b : _GEN_19653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19655 = 9'h113 == r_count_48_io_out ? io_r_275_b : _GEN_19654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19656 = 9'h114 == r_count_48_io_out ? io_r_276_b : _GEN_19655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19657 = 9'h115 == r_count_48_io_out ? io_r_277_b : _GEN_19656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19658 = 9'h116 == r_count_48_io_out ? io_r_278_b : _GEN_19657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19659 = 9'h117 == r_count_48_io_out ? io_r_279_b : _GEN_19658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19660 = 9'h118 == r_count_48_io_out ? io_r_280_b : _GEN_19659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19661 = 9'h119 == r_count_48_io_out ? io_r_281_b : _GEN_19660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19662 = 9'h11a == r_count_48_io_out ? io_r_282_b : _GEN_19661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19663 = 9'h11b == r_count_48_io_out ? io_r_283_b : _GEN_19662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19664 = 9'h11c == r_count_48_io_out ? io_r_284_b : _GEN_19663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19665 = 9'h11d == r_count_48_io_out ? io_r_285_b : _GEN_19664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19666 = 9'h11e == r_count_48_io_out ? io_r_286_b : _GEN_19665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19667 = 9'h11f == r_count_48_io_out ? io_r_287_b : _GEN_19666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19668 = 9'h120 == r_count_48_io_out ? io_r_288_b : _GEN_19667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19669 = 9'h121 == r_count_48_io_out ? io_r_289_b : _GEN_19668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19670 = 9'h122 == r_count_48_io_out ? io_r_290_b : _GEN_19669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19671 = 9'h123 == r_count_48_io_out ? io_r_291_b : _GEN_19670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19672 = 9'h124 == r_count_48_io_out ? io_r_292_b : _GEN_19671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19673 = 9'h125 == r_count_48_io_out ? io_r_293_b : _GEN_19672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19674 = 9'h126 == r_count_48_io_out ? io_r_294_b : _GEN_19673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19675 = 9'h127 == r_count_48_io_out ? io_r_295_b : _GEN_19674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19676 = 9'h128 == r_count_48_io_out ? io_r_296_b : _GEN_19675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19677 = 9'h129 == r_count_48_io_out ? io_r_297_b : _GEN_19676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19678 = 9'h12a == r_count_48_io_out ? io_r_298_b : _GEN_19677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19679 = 9'h12b == r_count_48_io_out ? io_r_299_b : _GEN_19678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19680 = 9'h12c == r_count_48_io_out ? io_r_300_b : _GEN_19679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19681 = 9'h12d == r_count_48_io_out ? io_r_301_b : _GEN_19680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19682 = 9'h12e == r_count_48_io_out ? io_r_302_b : _GEN_19681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19683 = 9'h12f == r_count_48_io_out ? io_r_303_b : _GEN_19682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19684 = 9'h130 == r_count_48_io_out ? io_r_304_b : _GEN_19683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19685 = 9'h131 == r_count_48_io_out ? io_r_305_b : _GEN_19684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19686 = 9'h132 == r_count_48_io_out ? io_r_306_b : _GEN_19685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19687 = 9'h133 == r_count_48_io_out ? io_r_307_b : _GEN_19686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19688 = 9'h134 == r_count_48_io_out ? io_r_308_b : _GEN_19687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19689 = 9'h135 == r_count_48_io_out ? io_r_309_b : _GEN_19688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19690 = 9'h136 == r_count_48_io_out ? io_r_310_b : _GEN_19689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19691 = 9'h137 == r_count_48_io_out ? io_r_311_b : _GEN_19690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19692 = 9'h138 == r_count_48_io_out ? io_r_312_b : _GEN_19691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19693 = 9'h139 == r_count_48_io_out ? io_r_313_b : _GEN_19692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19694 = 9'h13a == r_count_48_io_out ? io_r_314_b : _GEN_19693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19695 = 9'h13b == r_count_48_io_out ? io_r_315_b : _GEN_19694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19696 = 9'h13c == r_count_48_io_out ? io_r_316_b : _GEN_19695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19697 = 9'h13d == r_count_48_io_out ? io_r_317_b : _GEN_19696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19698 = 9'h13e == r_count_48_io_out ? io_r_318_b : _GEN_19697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19699 = 9'h13f == r_count_48_io_out ? io_r_319_b : _GEN_19698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19700 = 9'h140 == r_count_48_io_out ? io_r_320_b : _GEN_19699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19701 = 9'h141 == r_count_48_io_out ? io_r_321_b : _GEN_19700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19702 = 9'h142 == r_count_48_io_out ? io_r_322_b : _GEN_19701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19703 = 9'h143 == r_count_48_io_out ? io_r_323_b : _GEN_19702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19704 = 9'h144 == r_count_48_io_out ? io_r_324_b : _GEN_19703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19705 = 9'h145 == r_count_48_io_out ? io_r_325_b : _GEN_19704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19706 = 9'h146 == r_count_48_io_out ? io_r_326_b : _GEN_19705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19707 = 9'h147 == r_count_48_io_out ? io_r_327_b : _GEN_19706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19708 = 9'h148 == r_count_48_io_out ? io_r_328_b : _GEN_19707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19709 = 9'h149 == r_count_48_io_out ? io_r_329_b : _GEN_19708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19710 = 9'h14a == r_count_48_io_out ? io_r_330_b : _GEN_19709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19711 = 9'h14b == r_count_48_io_out ? io_r_331_b : _GEN_19710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19712 = 9'h14c == r_count_48_io_out ? io_r_332_b : _GEN_19711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19713 = 9'h14d == r_count_48_io_out ? io_r_333_b : _GEN_19712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19714 = 9'h14e == r_count_48_io_out ? io_r_334_b : _GEN_19713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19715 = 9'h14f == r_count_48_io_out ? io_r_335_b : _GEN_19714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19716 = 9'h150 == r_count_48_io_out ? io_r_336_b : _GEN_19715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19717 = 9'h151 == r_count_48_io_out ? io_r_337_b : _GEN_19716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19718 = 9'h152 == r_count_48_io_out ? io_r_338_b : _GEN_19717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19719 = 9'h153 == r_count_48_io_out ? io_r_339_b : _GEN_19718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19720 = 9'h154 == r_count_48_io_out ? io_r_340_b : _GEN_19719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19721 = 9'h155 == r_count_48_io_out ? io_r_341_b : _GEN_19720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19722 = 9'h156 == r_count_48_io_out ? io_r_342_b : _GEN_19721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19723 = 9'h157 == r_count_48_io_out ? io_r_343_b : _GEN_19722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19724 = 9'h158 == r_count_48_io_out ? io_r_344_b : _GEN_19723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19725 = 9'h159 == r_count_48_io_out ? io_r_345_b : _GEN_19724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19726 = 9'h15a == r_count_48_io_out ? io_r_346_b : _GEN_19725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19727 = 9'h15b == r_count_48_io_out ? io_r_347_b : _GEN_19726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19728 = 9'h15c == r_count_48_io_out ? io_r_348_b : _GEN_19727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19729 = 9'h15d == r_count_48_io_out ? io_r_349_b : _GEN_19728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19730 = 9'h15e == r_count_48_io_out ? io_r_350_b : _GEN_19729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19731 = 9'h15f == r_count_48_io_out ? io_r_351_b : _GEN_19730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19732 = 9'h160 == r_count_48_io_out ? io_r_352_b : _GEN_19731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19733 = 9'h161 == r_count_48_io_out ? io_r_353_b : _GEN_19732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19734 = 9'h162 == r_count_48_io_out ? io_r_354_b : _GEN_19733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19735 = 9'h163 == r_count_48_io_out ? io_r_355_b : _GEN_19734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19736 = 9'h164 == r_count_48_io_out ? io_r_356_b : _GEN_19735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19737 = 9'h165 == r_count_48_io_out ? io_r_357_b : _GEN_19736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19738 = 9'h166 == r_count_48_io_out ? io_r_358_b : _GEN_19737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19739 = 9'h167 == r_count_48_io_out ? io_r_359_b : _GEN_19738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19740 = 9'h168 == r_count_48_io_out ? io_r_360_b : _GEN_19739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19741 = 9'h169 == r_count_48_io_out ? io_r_361_b : _GEN_19740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19742 = 9'h16a == r_count_48_io_out ? io_r_362_b : _GEN_19741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19743 = 9'h16b == r_count_48_io_out ? io_r_363_b : _GEN_19742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19744 = 9'h16c == r_count_48_io_out ? io_r_364_b : _GEN_19743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19745 = 9'h16d == r_count_48_io_out ? io_r_365_b : _GEN_19744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19746 = 9'h16e == r_count_48_io_out ? io_r_366_b : _GEN_19745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19747 = 9'h16f == r_count_48_io_out ? io_r_367_b : _GEN_19746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19748 = 9'h170 == r_count_48_io_out ? io_r_368_b : _GEN_19747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19749 = 9'h171 == r_count_48_io_out ? io_r_369_b : _GEN_19748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19750 = 9'h172 == r_count_48_io_out ? io_r_370_b : _GEN_19749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19751 = 9'h173 == r_count_48_io_out ? io_r_371_b : _GEN_19750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19752 = 9'h174 == r_count_48_io_out ? io_r_372_b : _GEN_19751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19753 = 9'h175 == r_count_48_io_out ? io_r_373_b : _GEN_19752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19754 = 9'h176 == r_count_48_io_out ? io_r_374_b : _GEN_19753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19755 = 9'h177 == r_count_48_io_out ? io_r_375_b : _GEN_19754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19756 = 9'h178 == r_count_48_io_out ? io_r_376_b : _GEN_19755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19757 = 9'h179 == r_count_48_io_out ? io_r_377_b : _GEN_19756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19758 = 9'h17a == r_count_48_io_out ? io_r_378_b : _GEN_19757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19759 = 9'h17b == r_count_48_io_out ? io_r_379_b : _GEN_19758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19760 = 9'h17c == r_count_48_io_out ? io_r_380_b : _GEN_19759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19761 = 9'h17d == r_count_48_io_out ? io_r_381_b : _GEN_19760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19762 = 9'h17e == r_count_48_io_out ? io_r_382_b : _GEN_19761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19763 = 9'h17f == r_count_48_io_out ? io_r_383_b : _GEN_19762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19764 = 9'h180 == r_count_48_io_out ? io_r_384_b : _GEN_19763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19765 = 9'h181 == r_count_48_io_out ? io_r_385_b : _GEN_19764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19766 = 9'h182 == r_count_48_io_out ? io_r_386_b : _GEN_19765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19767 = 9'h183 == r_count_48_io_out ? io_r_387_b : _GEN_19766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19768 = 9'h184 == r_count_48_io_out ? io_r_388_b : _GEN_19767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19769 = 9'h185 == r_count_48_io_out ? io_r_389_b : _GEN_19768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19770 = 9'h186 == r_count_48_io_out ? io_r_390_b : _GEN_19769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19771 = 9'h187 == r_count_48_io_out ? io_r_391_b : _GEN_19770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19772 = 9'h188 == r_count_48_io_out ? io_r_392_b : _GEN_19771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19773 = 9'h189 == r_count_48_io_out ? io_r_393_b : _GEN_19772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19774 = 9'h18a == r_count_48_io_out ? io_r_394_b : _GEN_19773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19775 = 9'h18b == r_count_48_io_out ? io_r_395_b : _GEN_19774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19776 = 9'h18c == r_count_48_io_out ? io_r_396_b : _GEN_19775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19777 = 9'h18d == r_count_48_io_out ? io_r_397_b : _GEN_19776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19778 = 9'h18e == r_count_48_io_out ? io_r_398_b : _GEN_19777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19781 = 9'h1 == r_count_49_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19782 = 9'h2 == r_count_49_io_out ? io_r_2_b : _GEN_19781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19783 = 9'h3 == r_count_49_io_out ? io_r_3_b : _GEN_19782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19784 = 9'h4 == r_count_49_io_out ? io_r_4_b : _GEN_19783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19785 = 9'h5 == r_count_49_io_out ? io_r_5_b : _GEN_19784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19786 = 9'h6 == r_count_49_io_out ? io_r_6_b : _GEN_19785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19787 = 9'h7 == r_count_49_io_out ? io_r_7_b : _GEN_19786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19788 = 9'h8 == r_count_49_io_out ? io_r_8_b : _GEN_19787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19789 = 9'h9 == r_count_49_io_out ? io_r_9_b : _GEN_19788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19790 = 9'ha == r_count_49_io_out ? io_r_10_b : _GEN_19789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19791 = 9'hb == r_count_49_io_out ? io_r_11_b : _GEN_19790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19792 = 9'hc == r_count_49_io_out ? io_r_12_b : _GEN_19791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19793 = 9'hd == r_count_49_io_out ? io_r_13_b : _GEN_19792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19794 = 9'he == r_count_49_io_out ? io_r_14_b : _GEN_19793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19795 = 9'hf == r_count_49_io_out ? io_r_15_b : _GEN_19794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19796 = 9'h10 == r_count_49_io_out ? io_r_16_b : _GEN_19795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19797 = 9'h11 == r_count_49_io_out ? io_r_17_b : _GEN_19796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19798 = 9'h12 == r_count_49_io_out ? io_r_18_b : _GEN_19797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19799 = 9'h13 == r_count_49_io_out ? io_r_19_b : _GEN_19798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19800 = 9'h14 == r_count_49_io_out ? io_r_20_b : _GEN_19799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19801 = 9'h15 == r_count_49_io_out ? io_r_21_b : _GEN_19800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19802 = 9'h16 == r_count_49_io_out ? io_r_22_b : _GEN_19801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19803 = 9'h17 == r_count_49_io_out ? io_r_23_b : _GEN_19802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19804 = 9'h18 == r_count_49_io_out ? io_r_24_b : _GEN_19803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19805 = 9'h19 == r_count_49_io_out ? io_r_25_b : _GEN_19804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19806 = 9'h1a == r_count_49_io_out ? io_r_26_b : _GEN_19805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19807 = 9'h1b == r_count_49_io_out ? io_r_27_b : _GEN_19806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19808 = 9'h1c == r_count_49_io_out ? io_r_28_b : _GEN_19807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19809 = 9'h1d == r_count_49_io_out ? io_r_29_b : _GEN_19808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19810 = 9'h1e == r_count_49_io_out ? io_r_30_b : _GEN_19809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19811 = 9'h1f == r_count_49_io_out ? io_r_31_b : _GEN_19810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19812 = 9'h20 == r_count_49_io_out ? io_r_32_b : _GEN_19811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19813 = 9'h21 == r_count_49_io_out ? io_r_33_b : _GEN_19812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19814 = 9'h22 == r_count_49_io_out ? io_r_34_b : _GEN_19813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19815 = 9'h23 == r_count_49_io_out ? io_r_35_b : _GEN_19814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19816 = 9'h24 == r_count_49_io_out ? io_r_36_b : _GEN_19815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19817 = 9'h25 == r_count_49_io_out ? io_r_37_b : _GEN_19816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19818 = 9'h26 == r_count_49_io_out ? io_r_38_b : _GEN_19817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19819 = 9'h27 == r_count_49_io_out ? io_r_39_b : _GEN_19818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19820 = 9'h28 == r_count_49_io_out ? io_r_40_b : _GEN_19819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19821 = 9'h29 == r_count_49_io_out ? io_r_41_b : _GEN_19820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19822 = 9'h2a == r_count_49_io_out ? io_r_42_b : _GEN_19821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19823 = 9'h2b == r_count_49_io_out ? io_r_43_b : _GEN_19822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19824 = 9'h2c == r_count_49_io_out ? io_r_44_b : _GEN_19823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19825 = 9'h2d == r_count_49_io_out ? io_r_45_b : _GEN_19824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19826 = 9'h2e == r_count_49_io_out ? io_r_46_b : _GEN_19825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19827 = 9'h2f == r_count_49_io_out ? io_r_47_b : _GEN_19826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19828 = 9'h30 == r_count_49_io_out ? io_r_48_b : _GEN_19827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19829 = 9'h31 == r_count_49_io_out ? io_r_49_b : _GEN_19828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19830 = 9'h32 == r_count_49_io_out ? io_r_50_b : _GEN_19829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19831 = 9'h33 == r_count_49_io_out ? io_r_51_b : _GEN_19830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19832 = 9'h34 == r_count_49_io_out ? io_r_52_b : _GEN_19831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19833 = 9'h35 == r_count_49_io_out ? io_r_53_b : _GEN_19832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19834 = 9'h36 == r_count_49_io_out ? io_r_54_b : _GEN_19833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19835 = 9'h37 == r_count_49_io_out ? io_r_55_b : _GEN_19834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19836 = 9'h38 == r_count_49_io_out ? io_r_56_b : _GEN_19835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19837 = 9'h39 == r_count_49_io_out ? io_r_57_b : _GEN_19836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19838 = 9'h3a == r_count_49_io_out ? io_r_58_b : _GEN_19837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19839 = 9'h3b == r_count_49_io_out ? io_r_59_b : _GEN_19838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19840 = 9'h3c == r_count_49_io_out ? io_r_60_b : _GEN_19839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19841 = 9'h3d == r_count_49_io_out ? io_r_61_b : _GEN_19840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19842 = 9'h3e == r_count_49_io_out ? io_r_62_b : _GEN_19841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19843 = 9'h3f == r_count_49_io_out ? io_r_63_b : _GEN_19842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19844 = 9'h40 == r_count_49_io_out ? io_r_64_b : _GEN_19843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19845 = 9'h41 == r_count_49_io_out ? io_r_65_b : _GEN_19844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19846 = 9'h42 == r_count_49_io_out ? io_r_66_b : _GEN_19845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19847 = 9'h43 == r_count_49_io_out ? io_r_67_b : _GEN_19846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19848 = 9'h44 == r_count_49_io_out ? io_r_68_b : _GEN_19847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19849 = 9'h45 == r_count_49_io_out ? io_r_69_b : _GEN_19848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19850 = 9'h46 == r_count_49_io_out ? io_r_70_b : _GEN_19849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19851 = 9'h47 == r_count_49_io_out ? io_r_71_b : _GEN_19850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19852 = 9'h48 == r_count_49_io_out ? io_r_72_b : _GEN_19851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19853 = 9'h49 == r_count_49_io_out ? io_r_73_b : _GEN_19852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19854 = 9'h4a == r_count_49_io_out ? io_r_74_b : _GEN_19853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19855 = 9'h4b == r_count_49_io_out ? io_r_75_b : _GEN_19854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19856 = 9'h4c == r_count_49_io_out ? io_r_76_b : _GEN_19855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19857 = 9'h4d == r_count_49_io_out ? io_r_77_b : _GEN_19856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19858 = 9'h4e == r_count_49_io_out ? io_r_78_b : _GEN_19857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19859 = 9'h4f == r_count_49_io_out ? io_r_79_b : _GEN_19858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19860 = 9'h50 == r_count_49_io_out ? io_r_80_b : _GEN_19859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19861 = 9'h51 == r_count_49_io_out ? io_r_81_b : _GEN_19860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19862 = 9'h52 == r_count_49_io_out ? io_r_82_b : _GEN_19861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19863 = 9'h53 == r_count_49_io_out ? io_r_83_b : _GEN_19862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19864 = 9'h54 == r_count_49_io_out ? io_r_84_b : _GEN_19863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19865 = 9'h55 == r_count_49_io_out ? io_r_85_b : _GEN_19864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19866 = 9'h56 == r_count_49_io_out ? io_r_86_b : _GEN_19865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19867 = 9'h57 == r_count_49_io_out ? io_r_87_b : _GEN_19866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19868 = 9'h58 == r_count_49_io_out ? io_r_88_b : _GEN_19867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19869 = 9'h59 == r_count_49_io_out ? io_r_89_b : _GEN_19868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19870 = 9'h5a == r_count_49_io_out ? io_r_90_b : _GEN_19869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19871 = 9'h5b == r_count_49_io_out ? io_r_91_b : _GEN_19870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19872 = 9'h5c == r_count_49_io_out ? io_r_92_b : _GEN_19871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19873 = 9'h5d == r_count_49_io_out ? io_r_93_b : _GEN_19872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19874 = 9'h5e == r_count_49_io_out ? io_r_94_b : _GEN_19873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19875 = 9'h5f == r_count_49_io_out ? io_r_95_b : _GEN_19874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19876 = 9'h60 == r_count_49_io_out ? io_r_96_b : _GEN_19875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19877 = 9'h61 == r_count_49_io_out ? io_r_97_b : _GEN_19876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19878 = 9'h62 == r_count_49_io_out ? io_r_98_b : _GEN_19877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19879 = 9'h63 == r_count_49_io_out ? io_r_99_b : _GEN_19878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19880 = 9'h64 == r_count_49_io_out ? io_r_100_b : _GEN_19879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19881 = 9'h65 == r_count_49_io_out ? io_r_101_b : _GEN_19880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19882 = 9'h66 == r_count_49_io_out ? io_r_102_b : _GEN_19881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19883 = 9'h67 == r_count_49_io_out ? io_r_103_b : _GEN_19882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19884 = 9'h68 == r_count_49_io_out ? io_r_104_b : _GEN_19883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19885 = 9'h69 == r_count_49_io_out ? io_r_105_b : _GEN_19884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19886 = 9'h6a == r_count_49_io_out ? io_r_106_b : _GEN_19885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19887 = 9'h6b == r_count_49_io_out ? io_r_107_b : _GEN_19886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19888 = 9'h6c == r_count_49_io_out ? io_r_108_b : _GEN_19887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19889 = 9'h6d == r_count_49_io_out ? io_r_109_b : _GEN_19888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19890 = 9'h6e == r_count_49_io_out ? io_r_110_b : _GEN_19889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19891 = 9'h6f == r_count_49_io_out ? io_r_111_b : _GEN_19890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19892 = 9'h70 == r_count_49_io_out ? io_r_112_b : _GEN_19891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19893 = 9'h71 == r_count_49_io_out ? io_r_113_b : _GEN_19892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19894 = 9'h72 == r_count_49_io_out ? io_r_114_b : _GEN_19893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19895 = 9'h73 == r_count_49_io_out ? io_r_115_b : _GEN_19894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19896 = 9'h74 == r_count_49_io_out ? io_r_116_b : _GEN_19895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19897 = 9'h75 == r_count_49_io_out ? io_r_117_b : _GEN_19896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19898 = 9'h76 == r_count_49_io_out ? io_r_118_b : _GEN_19897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19899 = 9'h77 == r_count_49_io_out ? io_r_119_b : _GEN_19898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19900 = 9'h78 == r_count_49_io_out ? io_r_120_b : _GEN_19899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19901 = 9'h79 == r_count_49_io_out ? io_r_121_b : _GEN_19900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19902 = 9'h7a == r_count_49_io_out ? io_r_122_b : _GEN_19901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19903 = 9'h7b == r_count_49_io_out ? io_r_123_b : _GEN_19902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19904 = 9'h7c == r_count_49_io_out ? io_r_124_b : _GEN_19903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19905 = 9'h7d == r_count_49_io_out ? io_r_125_b : _GEN_19904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19906 = 9'h7e == r_count_49_io_out ? io_r_126_b : _GEN_19905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19907 = 9'h7f == r_count_49_io_out ? io_r_127_b : _GEN_19906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19908 = 9'h80 == r_count_49_io_out ? io_r_128_b : _GEN_19907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19909 = 9'h81 == r_count_49_io_out ? io_r_129_b : _GEN_19908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19910 = 9'h82 == r_count_49_io_out ? io_r_130_b : _GEN_19909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19911 = 9'h83 == r_count_49_io_out ? io_r_131_b : _GEN_19910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19912 = 9'h84 == r_count_49_io_out ? io_r_132_b : _GEN_19911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19913 = 9'h85 == r_count_49_io_out ? io_r_133_b : _GEN_19912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19914 = 9'h86 == r_count_49_io_out ? io_r_134_b : _GEN_19913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19915 = 9'h87 == r_count_49_io_out ? io_r_135_b : _GEN_19914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19916 = 9'h88 == r_count_49_io_out ? io_r_136_b : _GEN_19915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19917 = 9'h89 == r_count_49_io_out ? io_r_137_b : _GEN_19916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19918 = 9'h8a == r_count_49_io_out ? io_r_138_b : _GEN_19917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19919 = 9'h8b == r_count_49_io_out ? io_r_139_b : _GEN_19918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19920 = 9'h8c == r_count_49_io_out ? io_r_140_b : _GEN_19919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19921 = 9'h8d == r_count_49_io_out ? io_r_141_b : _GEN_19920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19922 = 9'h8e == r_count_49_io_out ? io_r_142_b : _GEN_19921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19923 = 9'h8f == r_count_49_io_out ? io_r_143_b : _GEN_19922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19924 = 9'h90 == r_count_49_io_out ? io_r_144_b : _GEN_19923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19925 = 9'h91 == r_count_49_io_out ? io_r_145_b : _GEN_19924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19926 = 9'h92 == r_count_49_io_out ? io_r_146_b : _GEN_19925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19927 = 9'h93 == r_count_49_io_out ? io_r_147_b : _GEN_19926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19928 = 9'h94 == r_count_49_io_out ? io_r_148_b : _GEN_19927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19929 = 9'h95 == r_count_49_io_out ? io_r_149_b : _GEN_19928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19930 = 9'h96 == r_count_49_io_out ? io_r_150_b : _GEN_19929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19931 = 9'h97 == r_count_49_io_out ? io_r_151_b : _GEN_19930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19932 = 9'h98 == r_count_49_io_out ? io_r_152_b : _GEN_19931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19933 = 9'h99 == r_count_49_io_out ? io_r_153_b : _GEN_19932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19934 = 9'h9a == r_count_49_io_out ? io_r_154_b : _GEN_19933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19935 = 9'h9b == r_count_49_io_out ? io_r_155_b : _GEN_19934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19936 = 9'h9c == r_count_49_io_out ? io_r_156_b : _GEN_19935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19937 = 9'h9d == r_count_49_io_out ? io_r_157_b : _GEN_19936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19938 = 9'h9e == r_count_49_io_out ? io_r_158_b : _GEN_19937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19939 = 9'h9f == r_count_49_io_out ? io_r_159_b : _GEN_19938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19940 = 9'ha0 == r_count_49_io_out ? io_r_160_b : _GEN_19939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19941 = 9'ha1 == r_count_49_io_out ? io_r_161_b : _GEN_19940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19942 = 9'ha2 == r_count_49_io_out ? io_r_162_b : _GEN_19941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19943 = 9'ha3 == r_count_49_io_out ? io_r_163_b : _GEN_19942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19944 = 9'ha4 == r_count_49_io_out ? io_r_164_b : _GEN_19943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19945 = 9'ha5 == r_count_49_io_out ? io_r_165_b : _GEN_19944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19946 = 9'ha6 == r_count_49_io_out ? io_r_166_b : _GEN_19945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19947 = 9'ha7 == r_count_49_io_out ? io_r_167_b : _GEN_19946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19948 = 9'ha8 == r_count_49_io_out ? io_r_168_b : _GEN_19947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19949 = 9'ha9 == r_count_49_io_out ? io_r_169_b : _GEN_19948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19950 = 9'haa == r_count_49_io_out ? io_r_170_b : _GEN_19949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19951 = 9'hab == r_count_49_io_out ? io_r_171_b : _GEN_19950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19952 = 9'hac == r_count_49_io_out ? io_r_172_b : _GEN_19951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19953 = 9'had == r_count_49_io_out ? io_r_173_b : _GEN_19952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19954 = 9'hae == r_count_49_io_out ? io_r_174_b : _GEN_19953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19955 = 9'haf == r_count_49_io_out ? io_r_175_b : _GEN_19954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19956 = 9'hb0 == r_count_49_io_out ? io_r_176_b : _GEN_19955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19957 = 9'hb1 == r_count_49_io_out ? io_r_177_b : _GEN_19956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19958 = 9'hb2 == r_count_49_io_out ? io_r_178_b : _GEN_19957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19959 = 9'hb3 == r_count_49_io_out ? io_r_179_b : _GEN_19958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19960 = 9'hb4 == r_count_49_io_out ? io_r_180_b : _GEN_19959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19961 = 9'hb5 == r_count_49_io_out ? io_r_181_b : _GEN_19960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19962 = 9'hb6 == r_count_49_io_out ? io_r_182_b : _GEN_19961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19963 = 9'hb7 == r_count_49_io_out ? io_r_183_b : _GEN_19962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19964 = 9'hb8 == r_count_49_io_out ? io_r_184_b : _GEN_19963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19965 = 9'hb9 == r_count_49_io_out ? io_r_185_b : _GEN_19964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19966 = 9'hba == r_count_49_io_out ? io_r_186_b : _GEN_19965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19967 = 9'hbb == r_count_49_io_out ? io_r_187_b : _GEN_19966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19968 = 9'hbc == r_count_49_io_out ? io_r_188_b : _GEN_19967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19969 = 9'hbd == r_count_49_io_out ? io_r_189_b : _GEN_19968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19970 = 9'hbe == r_count_49_io_out ? io_r_190_b : _GEN_19969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19971 = 9'hbf == r_count_49_io_out ? io_r_191_b : _GEN_19970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19972 = 9'hc0 == r_count_49_io_out ? io_r_192_b : _GEN_19971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19973 = 9'hc1 == r_count_49_io_out ? io_r_193_b : _GEN_19972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19974 = 9'hc2 == r_count_49_io_out ? io_r_194_b : _GEN_19973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19975 = 9'hc3 == r_count_49_io_out ? io_r_195_b : _GEN_19974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19976 = 9'hc4 == r_count_49_io_out ? io_r_196_b : _GEN_19975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19977 = 9'hc5 == r_count_49_io_out ? io_r_197_b : _GEN_19976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19978 = 9'hc6 == r_count_49_io_out ? io_r_198_b : _GEN_19977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19979 = 9'hc7 == r_count_49_io_out ? io_r_199_b : _GEN_19978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19980 = 9'hc8 == r_count_49_io_out ? io_r_200_b : _GEN_19979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19981 = 9'hc9 == r_count_49_io_out ? io_r_201_b : _GEN_19980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19982 = 9'hca == r_count_49_io_out ? io_r_202_b : _GEN_19981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19983 = 9'hcb == r_count_49_io_out ? io_r_203_b : _GEN_19982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19984 = 9'hcc == r_count_49_io_out ? io_r_204_b : _GEN_19983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19985 = 9'hcd == r_count_49_io_out ? io_r_205_b : _GEN_19984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19986 = 9'hce == r_count_49_io_out ? io_r_206_b : _GEN_19985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19987 = 9'hcf == r_count_49_io_out ? io_r_207_b : _GEN_19986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19988 = 9'hd0 == r_count_49_io_out ? io_r_208_b : _GEN_19987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19989 = 9'hd1 == r_count_49_io_out ? io_r_209_b : _GEN_19988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19990 = 9'hd2 == r_count_49_io_out ? io_r_210_b : _GEN_19989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19991 = 9'hd3 == r_count_49_io_out ? io_r_211_b : _GEN_19990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19992 = 9'hd4 == r_count_49_io_out ? io_r_212_b : _GEN_19991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19993 = 9'hd5 == r_count_49_io_out ? io_r_213_b : _GEN_19992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19994 = 9'hd6 == r_count_49_io_out ? io_r_214_b : _GEN_19993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19995 = 9'hd7 == r_count_49_io_out ? io_r_215_b : _GEN_19994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19996 = 9'hd8 == r_count_49_io_out ? io_r_216_b : _GEN_19995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19997 = 9'hd9 == r_count_49_io_out ? io_r_217_b : _GEN_19996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19998 = 9'hda == r_count_49_io_out ? io_r_218_b : _GEN_19997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19999 = 9'hdb == r_count_49_io_out ? io_r_219_b : _GEN_19998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20000 = 9'hdc == r_count_49_io_out ? io_r_220_b : _GEN_19999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20001 = 9'hdd == r_count_49_io_out ? io_r_221_b : _GEN_20000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20002 = 9'hde == r_count_49_io_out ? io_r_222_b : _GEN_20001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20003 = 9'hdf == r_count_49_io_out ? io_r_223_b : _GEN_20002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20004 = 9'he0 == r_count_49_io_out ? io_r_224_b : _GEN_20003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20005 = 9'he1 == r_count_49_io_out ? io_r_225_b : _GEN_20004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20006 = 9'he2 == r_count_49_io_out ? io_r_226_b : _GEN_20005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20007 = 9'he3 == r_count_49_io_out ? io_r_227_b : _GEN_20006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20008 = 9'he4 == r_count_49_io_out ? io_r_228_b : _GEN_20007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20009 = 9'he5 == r_count_49_io_out ? io_r_229_b : _GEN_20008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20010 = 9'he6 == r_count_49_io_out ? io_r_230_b : _GEN_20009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20011 = 9'he7 == r_count_49_io_out ? io_r_231_b : _GEN_20010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20012 = 9'he8 == r_count_49_io_out ? io_r_232_b : _GEN_20011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20013 = 9'he9 == r_count_49_io_out ? io_r_233_b : _GEN_20012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20014 = 9'hea == r_count_49_io_out ? io_r_234_b : _GEN_20013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20015 = 9'heb == r_count_49_io_out ? io_r_235_b : _GEN_20014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20016 = 9'hec == r_count_49_io_out ? io_r_236_b : _GEN_20015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20017 = 9'hed == r_count_49_io_out ? io_r_237_b : _GEN_20016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20018 = 9'hee == r_count_49_io_out ? io_r_238_b : _GEN_20017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20019 = 9'hef == r_count_49_io_out ? io_r_239_b : _GEN_20018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20020 = 9'hf0 == r_count_49_io_out ? io_r_240_b : _GEN_20019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20021 = 9'hf1 == r_count_49_io_out ? io_r_241_b : _GEN_20020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20022 = 9'hf2 == r_count_49_io_out ? io_r_242_b : _GEN_20021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20023 = 9'hf3 == r_count_49_io_out ? io_r_243_b : _GEN_20022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20024 = 9'hf4 == r_count_49_io_out ? io_r_244_b : _GEN_20023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20025 = 9'hf5 == r_count_49_io_out ? io_r_245_b : _GEN_20024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20026 = 9'hf6 == r_count_49_io_out ? io_r_246_b : _GEN_20025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20027 = 9'hf7 == r_count_49_io_out ? io_r_247_b : _GEN_20026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20028 = 9'hf8 == r_count_49_io_out ? io_r_248_b : _GEN_20027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20029 = 9'hf9 == r_count_49_io_out ? io_r_249_b : _GEN_20028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20030 = 9'hfa == r_count_49_io_out ? io_r_250_b : _GEN_20029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20031 = 9'hfb == r_count_49_io_out ? io_r_251_b : _GEN_20030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20032 = 9'hfc == r_count_49_io_out ? io_r_252_b : _GEN_20031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20033 = 9'hfd == r_count_49_io_out ? io_r_253_b : _GEN_20032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20034 = 9'hfe == r_count_49_io_out ? io_r_254_b : _GEN_20033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20035 = 9'hff == r_count_49_io_out ? io_r_255_b : _GEN_20034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20036 = 9'h100 == r_count_49_io_out ? io_r_256_b : _GEN_20035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20037 = 9'h101 == r_count_49_io_out ? io_r_257_b : _GEN_20036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20038 = 9'h102 == r_count_49_io_out ? io_r_258_b : _GEN_20037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20039 = 9'h103 == r_count_49_io_out ? io_r_259_b : _GEN_20038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20040 = 9'h104 == r_count_49_io_out ? io_r_260_b : _GEN_20039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20041 = 9'h105 == r_count_49_io_out ? io_r_261_b : _GEN_20040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20042 = 9'h106 == r_count_49_io_out ? io_r_262_b : _GEN_20041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20043 = 9'h107 == r_count_49_io_out ? io_r_263_b : _GEN_20042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20044 = 9'h108 == r_count_49_io_out ? io_r_264_b : _GEN_20043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20045 = 9'h109 == r_count_49_io_out ? io_r_265_b : _GEN_20044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20046 = 9'h10a == r_count_49_io_out ? io_r_266_b : _GEN_20045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20047 = 9'h10b == r_count_49_io_out ? io_r_267_b : _GEN_20046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20048 = 9'h10c == r_count_49_io_out ? io_r_268_b : _GEN_20047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20049 = 9'h10d == r_count_49_io_out ? io_r_269_b : _GEN_20048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20050 = 9'h10e == r_count_49_io_out ? io_r_270_b : _GEN_20049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20051 = 9'h10f == r_count_49_io_out ? io_r_271_b : _GEN_20050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20052 = 9'h110 == r_count_49_io_out ? io_r_272_b : _GEN_20051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20053 = 9'h111 == r_count_49_io_out ? io_r_273_b : _GEN_20052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20054 = 9'h112 == r_count_49_io_out ? io_r_274_b : _GEN_20053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20055 = 9'h113 == r_count_49_io_out ? io_r_275_b : _GEN_20054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20056 = 9'h114 == r_count_49_io_out ? io_r_276_b : _GEN_20055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20057 = 9'h115 == r_count_49_io_out ? io_r_277_b : _GEN_20056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20058 = 9'h116 == r_count_49_io_out ? io_r_278_b : _GEN_20057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20059 = 9'h117 == r_count_49_io_out ? io_r_279_b : _GEN_20058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20060 = 9'h118 == r_count_49_io_out ? io_r_280_b : _GEN_20059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20061 = 9'h119 == r_count_49_io_out ? io_r_281_b : _GEN_20060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20062 = 9'h11a == r_count_49_io_out ? io_r_282_b : _GEN_20061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20063 = 9'h11b == r_count_49_io_out ? io_r_283_b : _GEN_20062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20064 = 9'h11c == r_count_49_io_out ? io_r_284_b : _GEN_20063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20065 = 9'h11d == r_count_49_io_out ? io_r_285_b : _GEN_20064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20066 = 9'h11e == r_count_49_io_out ? io_r_286_b : _GEN_20065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20067 = 9'h11f == r_count_49_io_out ? io_r_287_b : _GEN_20066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20068 = 9'h120 == r_count_49_io_out ? io_r_288_b : _GEN_20067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20069 = 9'h121 == r_count_49_io_out ? io_r_289_b : _GEN_20068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20070 = 9'h122 == r_count_49_io_out ? io_r_290_b : _GEN_20069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20071 = 9'h123 == r_count_49_io_out ? io_r_291_b : _GEN_20070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20072 = 9'h124 == r_count_49_io_out ? io_r_292_b : _GEN_20071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20073 = 9'h125 == r_count_49_io_out ? io_r_293_b : _GEN_20072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20074 = 9'h126 == r_count_49_io_out ? io_r_294_b : _GEN_20073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20075 = 9'h127 == r_count_49_io_out ? io_r_295_b : _GEN_20074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20076 = 9'h128 == r_count_49_io_out ? io_r_296_b : _GEN_20075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20077 = 9'h129 == r_count_49_io_out ? io_r_297_b : _GEN_20076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20078 = 9'h12a == r_count_49_io_out ? io_r_298_b : _GEN_20077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20079 = 9'h12b == r_count_49_io_out ? io_r_299_b : _GEN_20078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20080 = 9'h12c == r_count_49_io_out ? io_r_300_b : _GEN_20079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20081 = 9'h12d == r_count_49_io_out ? io_r_301_b : _GEN_20080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20082 = 9'h12e == r_count_49_io_out ? io_r_302_b : _GEN_20081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20083 = 9'h12f == r_count_49_io_out ? io_r_303_b : _GEN_20082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20084 = 9'h130 == r_count_49_io_out ? io_r_304_b : _GEN_20083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20085 = 9'h131 == r_count_49_io_out ? io_r_305_b : _GEN_20084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20086 = 9'h132 == r_count_49_io_out ? io_r_306_b : _GEN_20085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20087 = 9'h133 == r_count_49_io_out ? io_r_307_b : _GEN_20086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20088 = 9'h134 == r_count_49_io_out ? io_r_308_b : _GEN_20087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20089 = 9'h135 == r_count_49_io_out ? io_r_309_b : _GEN_20088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20090 = 9'h136 == r_count_49_io_out ? io_r_310_b : _GEN_20089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20091 = 9'h137 == r_count_49_io_out ? io_r_311_b : _GEN_20090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20092 = 9'h138 == r_count_49_io_out ? io_r_312_b : _GEN_20091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20093 = 9'h139 == r_count_49_io_out ? io_r_313_b : _GEN_20092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20094 = 9'h13a == r_count_49_io_out ? io_r_314_b : _GEN_20093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20095 = 9'h13b == r_count_49_io_out ? io_r_315_b : _GEN_20094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20096 = 9'h13c == r_count_49_io_out ? io_r_316_b : _GEN_20095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20097 = 9'h13d == r_count_49_io_out ? io_r_317_b : _GEN_20096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20098 = 9'h13e == r_count_49_io_out ? io_r_318_b : _GEN_20097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20099 = 9'h13f == r_count_49_io_out ? io_r_319_b : _GEN_20098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20100 = 9'h140 == r_count_49_io_out ? io_r_320_b : _GEN_20099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20101 = 9'h141 == r_count_49_io_out ? io_r_321_b : _GEN_20100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20102 = 9'h142 == r_count_49_io_out ? io_r_322_b : _GEN_20101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20103 = 9'h143 == r_count_49_io_out ? io_r_323_b : _GEN_20102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20104 = 9'h144 == r_count_49_io_out ? io_r_324_b : _GEN_20103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20105 = 9'h145 == r_count_49_io_out ? io_r_325_b : _GEN_20104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20106 = 9'h146 == r_count_49_io_out ? io_r_326_b : _GEN_20105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20107 = 9'h147 == r_count_49_io_out ? io_r_327_b : _GEN_20106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20108 = 9'h148 == r_count_49_io_out ? io_r_328_b : _GEN_20107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20109 = 9'h149 == r_count_49_io_out ? io_r_329_b : _GEN_20108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20110 = 9'h14a == r_count_49_io_out ? io_r_330_b : _GEN_20109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20111 = 9'h14b == r_count_49_io_out ? io_r_331_b : _GEN_20110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20112 = 9'h14c == r_count_49_io_out ? io_r_332_b : _GEN_20111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20113 = 9'h14d == r_count_49_io_out ? io_r_333_b : _GEN_20112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20114 = 9'h14e == r_count_49_io_out ? io_r_334_b : _GEN_20113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20115 = 9'h14f == r_count_49_io_out ? io_r_335_b : _GEN_20114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20116 = 9'h150 == r_count_49_io_out ? io_r_336_b : _GEN_20115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20117 = 9'h151 == r_count_49_io_out ? io_r_337_b : _GEN_20116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20118 = 9'h152 == r_count_49_io_out ? io_r_338_b : _GEN_20117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20119 = 9'h153 == r_count_49_io_out ? io_r_339_b : _GEN_20118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20120 = 9'h154 == r_count_49_io_out ? io_r_340_b : _GEN_20119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20121 = 9'h155 == r_count_49_io_out ? io_r_341_b : _GEN_20120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20122 = 9'h156 == r_count_49_io_out ? io_r_342_b : _GEN_20121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20123 = 9'h157 == r_count_49_io_out ? io_r_343_b : _GEN_20122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20124 = 9'h158 == r_count_49_io_out ? io_r_344_b : _GEN_20123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20125 = 9'h159 == r_count_49_io_out ? io_r_345_b : _GEN_20124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20126 = 9'h15a == r_count_49_io_out ? io_r_346_b : _GEN_20125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20127 = 9'h15b == r_count_49_io_out ? io_r_347_b : _GEN_20126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20128 = 9'h15c == r_count_49_io_out ? io_r_348_b : _GEN_20127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20129 = 9'h15d == r_count_49_io_out ? io_r_349_b : _GEN_20128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20130 = 9'h15e == r_count_49_io_out ? io_r_350_b : _GEN_20129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20131 = 9'h15f == r_count_49_io_out ? io_r_351_b : _GEN_20130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20132 = 9'h160 == r_count_49_io_out ? io_r_352_b : _GEN_20131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20133 = 9'h161 == r_count_49_io_out ? io_r_353_b : _GEN_20132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20134 = 9'h162 == r_count_49_io_out ? io_r_354_b : _GEN_20133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20135 = 9'h163 == r_count_49_io_out ? io_r_355_b : _GEN_20134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20136 = 9'h164 == r_count_49_io_out ? io_r_356_b : _GEN_20135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20137 = 9'h165 == r_count_49_io_out ? io_r_357_b : _GEN_20136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20138 = 9'h166 == r_count_49_io_out ? io_r_358_b : _GEN_20137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20139 = 9'h167 == r_count_49_io_out ? io_r_359_b : _GEN_20138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20140 = 9'h168 == r_count_49_io_out ? io_r_360_b : _GEN_20139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20141 = 9'h169 == r_count_49_io_out ? io_r_361_b : _GEN_20140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20142 = 9'h16a == r_count_49_io_out ? io_r_362_b : _GEN_20141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20143 = 9'h16b == r_count_49_io_out ? io_r_363_b : _GEN_20142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20144 = 9'h16c == r_count_49_io_out ? io_r_364_b : _GEN_20143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20145 = 9'h16d == r_count_49_io_out ? io_r_365_b : _GEN_20144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20146 = 9'h16e == r_count_49_io_out ? io_r_366_b : _GEN_20145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20147 = 9'h16f == r_count_49_io_out ? io_r_367_b : _GEN_20146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20148 = 9'h170 == r_count_49_io_out ? io_r_368_b : _GEN_20147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20149 = 9'h171 == r_count_49_io_out ? io_r_369_b : _GEN_20148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20150 = 9'h172 == r_count_49_io_out ? io_r_370_b : _GEN_20149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20151 = 9'h173 == r_count_49_io_out ? io_r_371_b : _GEN_20150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20152 = 9'h174 == r_count_49_io_out ? io_r_372_b : _GEN_20151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20153 = 9'h175 == r_count_49_io_out ? io_r_373_b : _GEN_20152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20154 = 9'h176 == r_count_49_io_out ? io_r_374_b : _GEN_20153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20155 = 9'h177 == r_count_49_io_out ? io_r_375_b : _GEN_20154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20156 = 9'h178 == r_count_49_io_out ? io_r_376_b : _GEN_20155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20157 = 9'h179 == r_count_49_io_out ? io_r_377_b : _GEN_20156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20158 = 9'h17a == r_count_49_io_out ? io_r_378_b : _GEN_20157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20159 = 9'h17b == r_count_49_io_out ? io_r_379_b : _GEN_20158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20160 = 9'h17c == r_count_49_io_out ? io_r_380_b : _GEN_20159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20161 = 9'h17d == r_count_49_io_out ? io_r_381_b : _GEN_20160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20162 = 9'h17e == r_count_49_io_out ? io_r_382_b : _GEN_20161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20163 = 9'h17f == r_count_49_io_out ? io_r_383_b : _GEN_20162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20164 = 9'h180 == r_count_49_io_out ? io_r_384_b : _GEN_20163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20165 = 9'h181 == r_count_49_io_out ? io_r_385_b : _GEN_20164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20166 = 9'h182 == r_count_49_io_out ? io_r_386_b : _GEN_20165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20167 = 9'h183 == r_count_49_io_out ? io_r_387_b : _GEN_20166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20168 = 9'h184 == r_count_49_io_out ? io_r_388_b : _GEN_20167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20169 = 9'h185 == r_count_49_io_out ? io_r_389_b : _GEN_20168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20170 = 9'h186 == r_count_49_io_out ? io_r_390_b : _GEN_20169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20171 = 9'h187 == r_count_49_io_out ? io_r_391_b : _GEN_20170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20172 = 9'h188 == r_count_49_io_out ? io_r_392_b : _GEN_20171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20173 = 9'h189 == r_count_49_io_out ? io_r_393_b : _GEN_20172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20174 = 9'h18a == r_count_49_io_out ? io_r_394_b : _GEN_20173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20175 = 9'h18b == r_count_49_io_out ? io_r_395_b : _GEN_20174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20176 = 9'h18c == r_count_49_io_out ? io_r_396_b : _GEN_20175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20177 = 9'h18d == r_count_49_io_out ? io_r_397_b : _GEN_20176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20178 = 9'h18e == r_count_49_io_out ? io_r_398_b : _GEN_20177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20181 = 9'h1 == r_count_50_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20182 = 9'h2 == r_count_50_io_out ? io_r_2_b : _GEN_20181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20183 = 9'h3 == r_count_50_io_out ? io_r_3_b : _GEN_20182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20184 = 9'h4 == r_count_50_io_out ? io_r_4_b : _GEN_20183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20185 = 9'h5 == r_count_50_io_out ? io_r_5_b : _GEN_20184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20186 = 9'h6 == r_count_50_io_out ? io_r_6_b : _GEN_20185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20187 = 9'h7 == r_count_50_io_out ? io_r_7_b : _GEN_20186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20188 = 9'h8 == r_count_50_io_out ? io_r_8_b : _GEN_20187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20189 = 9'h9 == r_count_50_io_out ? io_r_9_b : _GEN_20188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20190 = 9'ha == r_count_50_io_out ? io_r_10_b : _GEN_20189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20191 = 9'hb == r_count_50_io_out ? io_r_11_b : _GEN_20190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20192 = 9'hc == r_count_50_io_out ? io_r_12_b : _GEN_20191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20193 = 9'hd == r_count_50_io_out ? io_r_13_b : _GEN_20192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20194 = 9'he == r_count_50_io_out ? io_r_14_b : _GEN_20193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20195 = 9'hf == r_count_50_io_out ? io_r_15_b : _GEN_20194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20196 = 9'h10 == r_count_50_io_out ? io_r_16_b : _GEN_20195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20197 = 9'h11 == r_count_50_io_out ? io_r_17_b : _GEN_20196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20198 = 9'h12 == r_count_50_io_out ? io_r_18_b : _GEN_20197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20199 = 9'h13 == r_count_50_io_out ? io_r_19_b : _GEN_20198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20200 = 9'h14 == r_count_50_io_out ? io_r_20_b : _GEN_20199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20201 = 9'h15 == r_count_50_io_out ? io_r_21_b : _GEN_20200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20202 = 9'h16 == r_count_50_io_out ? io_r_22_b : _GEN_20201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20203 = 9'h17 == r_count_50_io_out ? io_r_23_b : _GEN_20202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20204 = 9'h18 == r_count_50_io_out ? io_r_24_b : _GEN_20203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20205 = 9'h19 == r_count_50_io_out ? io_r_25_b : _GEN_20204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20206 = 9'h1a == r_count_50_io_out ? io_r_26_b : _GEN_20205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20207 = 9'h1b == r_count_50_io_out ? io_r_27_b : _GEN_20206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20208 = 9'h1c == r_count_50_io_out ? io_r_28_b : _GEN_20207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20209 = 9'h1d == r_count_50_io_out ? io_r_29_b : _GEN_20208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20210 = 9'h1e == r_count_50_io_out ? io_r_30_b : _GEN_20209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20211 = 9'h1f == r_count_50_io_out ? io_r_31_b : _GEN_20210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20212 = 9'h20 == r_count_50_io_out ? io_r_32_b : _GEN_20211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20213 = 9'h21 == r_count_50_io_out ? io_r_33_b : _GEN_20212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20214 = 9'h22 == r_count_50_io_out ? io_r_34_b : _GEN_20213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20215 = 9'h23 == r_count_50_io_out ? io_r_35_b : _GEN_20214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20216 = 9'h24 == r_count_50_io_out ? io_r_36_b : _GEN_20215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20217 = 9'h25 == r_count_50_io_out ? io_r_37_b : _GEN_20216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20218 = 9'h26 == r_count_50_io_out ? io_r_38_b : _GEN_20217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20219 = 9'h27 == r_count_50_io_out ? io_r_39_b : _GEN_20218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20220 = 9'h28 == r_count_50_io_out ? io_r_40_b : _GEN_20219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20221 = 9'h29 == r_count_50_io_out ? io_r_41_b : _GEN_20220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20222 = 9'h2a == r_count_50_io_out ? io_r_42_b : _GEN_20221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20223 = 9'h2b == r_count_50_io_out ? io_r_43_b : _GEN_20222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20224 = 9'h2c == r_count_50_io_out ? io_r_44_b : _GEN_20223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20225 = 9'h2d == r_count_50_io_out ? io_r_45_b : _GEN_20224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20226 = 9'h2e == r_count_50_io_out ? io_r_46_b : _GEN_20225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20227 = 9'h2f == r_count_50_io_out ? io_r_47_b : _GEN_20226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20228 = 9'h30 == r_count_50_io_out ? io_r_48_b : _GEN_20227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20229 = 9'h31 == r_count_50_io_out ? io_r_49_b : _GEN_20228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20230 = 9'h32 == r_count_50_io_out ? io_r_50_b : _GEN_20229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20231 = 9'h33 == r_count_50_io_out ? io_r_51_b : _GEN_20230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20232 = 9'h34 == r_count_50_io_out ? io_r_52_b : _GEN_20231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20233 = 9'h35 == r_count_50_io_out ? io_r_53_b : _GEN_20232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20234 = 9'h36 == r_count_50_io_out ? io_r_54_b : _GEN_20233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20235 = 9'h37 == r_count_50_io_out ? io_r_55_b : _GEN_20234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20236 = 9'h38 == r_count_50_io_out ? io_r_56_b : _GEN_20235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20237 = 9'h39 == r_count_50_io_out ? io_r_57_b : _GEN_20236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20238 = 9'h3a == r_count_50_io_out ? io_r_58_b : _GEN_20237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20239 = 9'h3b == r_count_50_io_out ? io_r_59_b : _GEN_20238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20240 = 9'h3c == r_count_50_io_out ? io_r_60_b : _GEN_20239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20241 = 9'h3d == r_count_50_io_out ? io_r_61_b : _GEN_20240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20242 = 9'h3e == r_count_50_io_out ? io_r_62_b : _GEN_20241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20243 = 9'h3f == r_count_50_io_out ? io_r_63_b : _GEN_20242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20244 = 9'h40 == r_count_50_io_out ? io_r_64_b : _GEN_20243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20245 = 9'h41 == r_count_50_io_out ? io_r_65_b : _GEN_20244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20246 = 9'h42 == r_count_50_io_out ? io_r_66_b : _GEN_20245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20247 = 9'h43 == r_count_50_io_out ? io_r_67_b : _GEN_20246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20248 = 9'h44 == r_count_50_io_out ? io_r_68_b : _GEN_20247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20249 = 9'h45 == r_count_50_io_out ? io_r_69_b : _GEN_20248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20250 = 9'h46 == r_count_50_io_out ? io_r_70_b : _GEN_20249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20251 = 9'h47 == r_count_50_io_out ? io_r_71_b : _GEN_20250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20252 = 9'h48 == r_count_50_io_out ? io_r_72_b : _GEN_20251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20253 = 9'h49 == r_count_50_io_out ? io_r_73_b : _GEN_20252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20254 = 9'h4a == r_count_50_io_out ? io_r_74_b : _GEN_20253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20255 = 9'h4b == r_count_50_io_out ? io_r_75_b : _GEN_20254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20256 = 9'h4c == r_count_50_io_out ? io_r_76_b : _GEN_20255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20257 = 9'h4d == r_count_50_io_out ? io_r_77_b : _GEN_20256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20258 = 9'h4e == r_count_50_io_out ? io_r_78_b : _GEN_20257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20259 = 9'h4f == r_count_50_io_out ? io_r_79_b : _GEN_20258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20260 = 9'h50 == r_count_50_io_out ? io_r_80_b : _GEN_20259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20261 = 9'h51 == r_count_50_io_out ? io_r_81_b : _GEN_20260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20262 = 9'h52 == r_count_50_io_out ? io_r_82_b : _GEN_20261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20263 = 9'h53 == r_count_50_io_out ? io_r_83_b : _GEN_20262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20264 = 9'h54 == r_count_50_io_out ? io_r_84_b : _GEN_20263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20265 = 9'h55 == r_count_50_io_out ? io_r_85_b : _GEN_20264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20266 = 9'h56 == r_count_50_io_out ? io_r_86_b : _GEN_20265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20267 = 9'h57 == r_count_50_io_out ? io_r_87_b : _GEN_20266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20268 = 9'h58 == r_count_50_io_out ? io_r_88_b : _GEN_20267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20269 = 9'h59 == r_count_50_io_out ? io_r_89_b : _GEN_20268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20270 = 9'h5a == r_count_50_io_out ? io_r_90_b : _GEN_20269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20271 = 9'h5b == r_count_50_io_out ? io_r_91_b : _GEN_20270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20272 = 9'h5c == r_count_50_io_out ? io_r_92_b : _GEN_20271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20273 = 9'h5d == r_count_50_io_out ? io_r_93_b : _GEN_20272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20274 = 9'h5e == r_count_50_io_out ? io_r_94_b : _GEN_20273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20275 = 9'h5f == r_count_50_io_out ? io_r_95_b : _GEN_20274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20276 = 9'h60 == r_count_50_io_out ? io_r_96_b : _GEN_20275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20277 = 9'h61 == r_count_50_io_out ? io_r_97_b : _GEN_20276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20278 = 9'h62 == r_count_50_io_out ? io_r_98_b : _GEN_20277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20279 = 9'h63 == r_count_50_io_out ? io_r_99_b : _GEN_20278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20280 = 9'h64 == r_count_50_io_out ? io_r_100_b : _GEN_20279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20281 = 9'h65 == r_count_50_io_out ? io_r_101_b : _GEN_20280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20282 = 9'h66 == r_count_50_io_out ? io_r_102_b : _GEN_20281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20283 = 9'h67 == r_count_50_io_out ? io_r_103_b : _GEN_20282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20284 = 9'h68 == r_count_50_io_out ? io_r_104_b : _GEN_20283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20285 = 9'h69 == r_count_50_io_out ? io_r_105_b : _GEN_20284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20286 = 9'h6a == r_count_50_io_out ? io_r_106_b : _GEN_20285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20287 = 9'h6b == r_count_50_io_out ? io_r_107_b : _GEN_20286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20288 = 9'h6c == r_count_50_io_out ? io_r_108_b : _GEN_20287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20289 = 9'h6d == r_count_50_io_out ? io_r_109_b : _GEN_20288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20290 = 9'h6e == r_count_50_io_out ? io_r_110_b : _GEN_20289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20291 = 9'h6f == r_count_50_io_out ? io_r_111_b : _GEN_20290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20292 = 9'h70 == r_count_50_io_out ? io_r_112_b : _GEN_20291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20293 = 9'h71 == r_count_50_io_out ? io_r_113_b : _GEN_20292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20294 = 9'h72 == r_count_50_io_out ? io_r_114_b : _GEN_20293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20295 = 9'h73 == r_count_50_io_out ? io_r_115_b : _GEN_20294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20296 = 9'h74 == r_count_50_io_out ? io_r_116_b : _GEN_20295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20297 = 9'h75 == r_count_50_io_out ? io_r_117_b : _GEN_20296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20298 = 9'h76 == r_count_50_io_out ? io_r_118_b : _GEN_20297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20299 = 9'h77 == r_count_50_io_out ? io_r_119_b : _GEN_20298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20300 = 9'h78 == r_count_50_io_out ? io_r_120_b : _GEN_20299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20301 = 9'h79 == r_count_50_io_out ? io_r_121_b : _GEN_20300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20302 = 9'h7a == r_count_50_io_out ? io_r_122_b : _GEN_20301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20303 = 9'h7b == r_count_50_io_out ? io_r_123_b : _GEN_20302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20304 = 9'h7c == r_count_50_io_out ? io_r_124_b : _GEN_20303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20305 = 9'h7d == r_count_50_io_out ? io_r_125_b : _GEN_20304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20306 = 9'h7e == r_count_50_io_out ? io_r_126_b : _GEN_20305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20307 = 9'h7f == r_count_50_io_out ? io_r_127_b : _GEN_20306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20308 = 9'h80 == r_count_50_io_out ? io_r_128_b : _GEN_20307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20309 = 9'h81 == r_count_50_io_out ? io_r_129_b : _GEN_20308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20310 = 9'h82 == r_count_50_io_out ? io_r_130_b : _GEN_20309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20311 = 9'h83 == r_count_50_io_out ? io_r_131_b : _GEN_20310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20312 = 9'h84 == r_count_50_io_out ? io_r_132_b : _GEN_20311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20313 = 9'h85 == r_count_50_io_out ? io_r_133_b : _GEN_20312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20314 = 9'h86 == r_count_50_io_out ? io_r_134_b : _GEN_20313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20315 = 9'h87 == r_count_50_io_out ? io_r_135_b : _GEN_20314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20316 = 9'h88 == r_count_50_io_out ? io_r_136_b : _GEN_20315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20317 = 9'h89 == r_count_50_io_out ? io_r_137_b : _GEN_20316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20318 = 9'h8a == r_count_50_io_out ? io_r_138_b : _GEN_20317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20319 = 9'h8b == r_count_50_io_out ? io_r_139_b : _GEN_20318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20320 = 9'h8c == r_count_50_io_out ? io_r_140_b : _GEN_20319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20321 = 9'h8d == r_count_50_io_out ? io_r_141_b : _GEN_20320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20322 = 9'h8e == r_count_50_io_out ? io_r_142_b : _GEN_20321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20323 = 9'h8f == r_count_50_io_out ? io_r_143_b : _GEN_20322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20324 = 9'h90 == r_count_50_io_out ? io_r_144_b : _GEN_20323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20325 = 9'h91 == r_count_50_io_out ? io_r_145_b : _GEN_20324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20326 = 9'h92 == r_count_50_io_out ? io_r_146_b : _GEN_20325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20327 = 9'h93 == r_count_50_io_out ? io_r_147_b : _GEN_20326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20328 = 9'h94 == r_count_50_io_out ? io_r_148_b : _GEN_20327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20329 = 9'h95 == r_count_50_io_out ? io_r_149_b : _GEN_20328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20330 = 9'h96 == r_count_50_io_out ? io_r_150_b : _GEN_20329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20331 = 9'h97 == r_count_50_io_out ? io_r_151_b : _GEN_20330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20332 = 9'h98 == r_count_50_io_out ? io_r_152_b : _GEN_20331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20333 = 9'h99 == r_count_50_io_out ? io_r_153_b : _GEN_20332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20334 = 9'h9a == r_count_50_io_out ? io_r_154_b : _GEN_20333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20335 = 9'h9b == r_count_50_io_out ? io_r_155_b : _GEN_20334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20336 = 9'h9c == r_count_50_io_out ? io_r_156_b : _GEN_20335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20337 = 9'h9d == r_count_50_io_out ? io_r_157_b : _GEN_20336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20338 = 9'h9e == r_count_50_io_out ? io_r_158_b : _GEN_20337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20339 = 9'h9f == r_count_50_io_out ? io_r_159_b : _GEN_20338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20340 = 9'ha0 == r_count_50_io_out ? io_r_160_b : _GEN_20339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20341 = 9'ha1 == r_count_50_io_out ? io_r_161_b : _GEN_20340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20342 = 9'ha2 == r_count_50_io_out ? io_r_162_b : _GEN_20341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20343 = 9'ha3 == r_count_50_io_out ? io_r_163_b : _GEN_20342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20344 = 9'ha4 == r_count_50_io_out ? io_r_164_b : _GEN_20343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20345 = 9'ha5 == r_count_50_io_out ? io_r_165_b : _GEN_20344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20346 = 9'ha6 == r_count_50_io_out ? io_r_166_b : _GEN_20345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20347 = 9'ha7 == r_count_50_io_out ? io_r_167_b : _GEN_20346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20348 = 9'ha8 == r_count_50_io_out ? io_r_168_b : _GEN_20347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20349 = 9'ha9 == r_count_50_io_out ? io_r_169_b : _GEN_20348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20350 = 9'haa == r_count_50_io_out ? io_r_170_b : _GEN_20349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20351 = 9'hab == r_count_50_io_out ? io_r_171_b : _GEN_20350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20352 = 9'hac == r_count_50_io_out ? io_r_172_b : _GEN_20351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20353 = 9'had == r_count_50_io_out ? io_r_173_b : _GEN_20352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20354 = 9'hae == r_count_50_io_out ? io_r_174_b : _GEN_20353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20355 = 9'haf == r_count_50_io_out ? io_r_175_b : _GEN_20354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20356 = 9'hb0 == r_count_50_io_out ? io_r_176_b : _GEN_20355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20357 = 9'hb1 == r_count_50_io_out ? io_r_177_b : _GEN_20356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20358 = 9'hb2 == r_count_50_io_out ? io_r_178_b : _GEN_20357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20359 = 9'hb3 == r_count_50_io_out ? io_r_179_b : _GEN_20358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20360 = 9'hb4 == r_count_50_io_out ? io_r_180_b : _GEN_20359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20361 = 9'hb5 == r_count_50_io_out ? io_r_181_b : _GEN_20360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20362 = 9'hb6 == r_count_50_io_out ? io_r_182_b : _GEN_20361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20363 = 9'hb7 == r_count_50_io_out ? io_r_183_b : _GEN_20362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20364 = 9'hb8 == r_count_50_io_out ? io_r_184_b : _GEN_20363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20365 = 9'hb9 == r_count_50_io_out ? io_r_185_b : _GEN_20364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20366 = 9'hba == r_count_50_io_out ? io_r_186_b : _GEN_20365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20367 = 9'hbb == r_count_50_io_out ? io_r_187_b : _GEN_20366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20368 = 9'hbc == r_count_50_io_out ? io_r_188_b : _GEN_20367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20369 = 9'hbd == r_count_50_io_out ? io_r_189_b : _GEN_20368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20370 = 9'hbe == r_count_50_io_out ? io_r_190_b : _GEN_20369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20371 = 9'hbf == r_count_50_io_out ? io_r_191_b : _GEN_20370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20372 = 9'hc0 == r_count_50_io_out ? io_r_192_b : _GEN_20371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20373 = 9'hc1 == r_count_50_io_out ? io_r_193_b : _GEN_20372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20374 = 9'hc2 == r_count_50_io_out ? io_r_194_b : _GEN_20373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20375 = 9'hc3 == r_count_50_io_out ? io_r_195_b : _GEN_20374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20376 = 9'hc4 == r_count_50_io_out ? io_r_196_b : _GEN_20375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20377 = 9'hc5 == r_count_50_io_out ? io_r_197_b : _GEN_20376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20378 = 9'hc6 == r_count_50_io_out ? io_r_198_b : _GEN_20377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20379 = 9'hc7 == r_count_50_io_out ? io_r_199_b : _GEN_20378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20380 = 9'hc8 == r_count_50_io_out ? io_r_200_b : _GEN_20379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20381 = 9'hc9 == r_count_50_io_out ? io_r_201_b : _GEN_20380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20382 = 9'hca == r_count_50_io_out ? io_r_202_b : _GEN_20381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20383 = 9'hcb == r_count_50_io_out ? io_r_203_b : _GEN_20382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20384 = 9'hcc == r_count_50_io_out ? io_r_204_b : _GEN_20383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20385 = 9'hcd == r_count_50_io_out ? io_r_205_b : _GEN_20384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20386 = 9'hce == r_count_50_io_out ? io_r_206_b : _GEN_20385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20387 = 9'hcf == r_count_50_io_out ? io_r_207_b : _GEN_20386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20388 = 9'hd0 == r_count_50_io_out ? io_r_208_b : _GEN_20387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20389 = 9'hd1 == r_count_50_io_out ? io_r_209_b : _GEN_20388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20390 = 9'hd2 == r_count_50_io_out ? io_r_210_b : _GEN_20389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20391 = 9'hd3 == r_count_50_io_out ? io_r_211_b : _GEN_20390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20392 = 9'hd4 == r_count_50_io_out ? io_r_212_b : _GEN_20391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20393 = 9'hd5 == r_count_50_io_out ? io_r_213_b : _GEN_20392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20394 = 9'hd6 == r_count_50_io_out ? io_r_214_b : _GEN_20393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20395 = 9'hd7 == r_count_50_io_out ? io_r_215_b : _GEN_20394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20396 = 9'hd8 == r_count_50_io_out ? io_r_216_b : _GEN_20395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20397 = 9'hd9 == r_count_50_io_out ? io_r_217_b : _GEN_20396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20398 = 9'hda == r_count_50_io_out ? io_r_218_b : _GEN_20397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20399 = 9'hdb == r_count_50_io_out ? io_r_219_b : _GEN_20398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20400 = 9'hdc == r_count_50_io_out ? io_r_220_b : _GEN_20399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20401 = 9'hdd == r_count_50_io_out ? io_r_221_b : _GEN_20400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20402 = 9'hde == r_count_50_io_out ? io_r_222_b : _GEN_20401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20403 = 9'hdf == r_count_50_io_out ? io_r_223_b : _GEN_20402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20404 = 9'he0 == r_count_50_io_out ? io_r_224_b : _GEN_20403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20405 = 9'he1 == r_count_50_io_out ? io_r_225_b : _GEN_20404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20406 = 9'he2 == r_count_50_io_out ? io_r_226_b : _GEN_20405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20407 = 9'he3 == r_count_50_io_out ? io_r_227_b : _GEN_20406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20408 = 9'he4 == r_count_50_io_out ? io_r_228_b : _GEN_20407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20409 = 9'he5 == r_count_50_io_out ? io_r_229_b : _GEN_20408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20410 = 9'he6 == r_count_50_io_out ? io_r_230_b : _GEN_20409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20411 = 9'he7 == r_count_50_io_out ? io_r_231_b : _GEN_20410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20412 = 9'he8 == r_count_50_io_out ? io_r_232_b : _GEN_20411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20413 = 9'he9 == r_count_50_io_out ? io_r_233_b : _GEN_20412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20414 = 9'hea == r_count_50_io_out ? io_r_234_b : _GEN_20413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20415 = 9'heb == r_count_50_io_out ? io_r_235_b : _GEN_20414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20416 = 9'hec == r_count_50_io_out ? io_r_236_b : _GEN_20415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20417 = 9'hed == r_count_50_io_out ? io_r_237_b : _GEN_20416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20418 = 9'hee == r_count_50_io_out ? io_r_238_b : _GEN_20417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20419 = 9'hef == r_count_50_io_out ? io_r_239_b : _GEN_20418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20420 = 9'hf0 == r_count_50_io_out ? io_r_240_b : _GEN_20419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20421 = 9'hf1 == r_count_50_io_out ? io_r_241_b : _GEN_20420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20422 = 9'hf2 == r_count_50_io_out ? io_r_242_b : _GEN_20421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20423 = 9'hf3 == r_count_50_io_out ? io_r_243_b : _GEN_20422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20424 = 9'hf4 == r_count_50_io_out ? io_r_244_b : _GEN_20423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20425 = 9'hf5 == r_count_50_io_out ? io_r_245_b : _GEN_20424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20426 = 9'hf6 == r_count_50_io_out ? io_r_246_b : _GEN_20425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20427 = 9'hf7 == r_count_50_io_out ? io_r_247_b : _GEN_20426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20428 = 9'hf8 == r_count_50_io_out ? io_r_248_b : _GEN_20427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20429 = 9'hf9 == r_count_50_io_out ? io_r_249_b : _GEN_20428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20430 = 9'hfa == r_count_50_io_out ? io_r_250_b : _GEN_20429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20431 = 9'hfb == r_count_50_io_out ? io_r_251_b : _GEN_20430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20432 = 9'hfc == r_count_50_io_out ? io_r_252_b : _GEN_20431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20433 = 9'hfd == r_count_50_io_out ? io_r_253_b : _GEN_20432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20434 = 9'hfe == r_count_50_io_out ? io_r_254_b : _GEN_20433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20435 = 9'hff == r_count_50_io_out ? io_r_255_b : _GEN_20434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20436 = 9'h100 == r_count_50_io_out ? io_r_256_b : _GEN_20435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20437 = 9'h101 == r_count_50_io_out ? io_r_257_b : _GEN_20436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20438 = 9'h102 == r_count_50_io_out ? io_r_258_b : _GEN_20437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20439 = 9'h103 == r_count_50_io_out ? io_r_259_b : _GEN_20438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20440 = 9'h104 == r_count_50_io_out ? io_r_260_b : _GEN_20439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20441 = 9'h105 == r_count_50_io_out ? io_r_261_b : _GEN_20440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20442 = 9'h106 == r_count_50_io_out ? io_r_262_b : _GEN_20441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20443 = 9'h107 == r_count_50_io_out ? io_r_263_b : _GEN_20442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20444 = 9'h108 == r_count_50_io_out ? io_r_264_b : _GEN_20443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20445 = 9'h109 == r_count_50_io_out ? io_r_265_b : _GEN_20444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20446 = 9'h10a == r_count_50_io_out ? io_r_266_b : _GEN_20445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20447 = 9'h10b == r_count_50_io_out ? io_r_267_b : _GEN_20446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20448 = 9'h10c == r_count_50_io_out ? io_r_268_b : _GEN_20447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20449 = 9'h10d == r_count_50_io_out ? io_r_269_b : _GEN_20448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20450 = 9'h10e == r_count_50_io_out ? io_r_270_b : _GEN_20449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20451 = 9'h10f == r_count_50_io_out ? io_r_271_b : _GEN_20450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20452 = 9'h110 == r_count_50_io_out ? io_r_272_b : _GEN_20451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20453 = 9'h111 == r_count_50_io_out ? io_r_273_b : _GEN_20452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20454 = 9'h112 == r_count_50_io_out ? io_r_274_b : _GEN_20453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20455 = 9'h113 == r_count_50_io_out ? io_r_275_b : _GEN_20454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20456 = 9'h114 == r_count_50_io_out ? io_r_276_b : _GEN_20455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20457 = 9'h115 == r_count_50_io_out ? io_r_277_b : _GEN_20456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20458 = 9'h116 == r_count_50_io_out ? io_r_278_b : _GEN_20457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20459 = 9'h117 == r_count_50_io_out ? io_r_279_b : _GEN_20458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20460 = 9'h118 == r_count_50_io_out ? io_r_280_b : _GEN_20459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20461 = 9'h119 == r_count_50_io_out ? io_r_281_b : _GEN_20460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20462 = 9'h11a == r_count_50_io_out ? io_r_282_b : _GEN_20461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20463 = 9'h11b == r_count_50_io_out ? io_r_283_b : _GEN_20462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20464 = 9'h11c == r_count_50_io_out ? io_r_284_b : _GEN_20463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20465 = 9'h11d == r_count_50_io_out ? io_r_285_b : _GEN_20464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20466 = 9'h11e == r_count_50_io_out ? io_r_286_b : _GEN_20465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20467 = 9'h11f == r_count_50_io_out ? io_r_287_b : _GEN_20466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20468 = 9'h120 == r_count_50_io_out ? io_r_288_b : _GEN_20467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20469 = 9'h121 == r_count_50_io_out ? io_r_289_b : _GEN_20468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20470 = 9'h122 == r_count_50_io_out ? io_r_290_b : _GEN_20469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20471 = 9'h123 == r_count_50_io_out ? io_r_291_b : _GEN_20470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20472 = 9'h124 == r_count_50_io_out ? io_r_292_b : _GEN_20471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20473 = 9'h125 == r_count_50_io_out ? io_r_293_b : _GEN_20472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20474 = 9'h126 == r_count_50_io_out ? io_r_294_b : _GEN_20473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20475 = 9'h127 == r_count_50_io_out ? io_r_295_b : _GEN_20474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20476 = 9'h128 == r_count_50_io_out ? io_r_296_b : _GEN_20475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20477 = 9'h129 == r_count_50_io_out ? io_r_297_b : _GEN_20476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20478 = 9'h12a == r_count_50_io_out ? io_r_298_b : _GEN_20477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20479 = 9'h12b == r_count_50_io_out ? io_r_299_b : _GEN_20478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20480 = 9'h12c == r_count_50_io_out ? io_r_300_b : _GEN_20479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20481 = 9'h12d == r_count_50_io_out ? io_r_301_b : _GEN_20480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20482 = 9'h12e == r_count_50_io_out ? io_r_302_b : _GEN_20481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20483 = 9'h12f == r_count_50_io_out ? io_r_303_b : _GEN_20482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20484 = 9'h130 == r_count_50_io_out ? io_r_304_b : _GEN_20483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20485 = 9'h131 == r_count_50_io_out ? io_r_305_b : _GEN_20484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20486 = 9'h132 == r_count_50_io_out ? io_r_306_b : _GEN_20485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20487 = 9'h133 == r_count_50_io_out ? io_r_307_b : _GEN_20486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20488 = 9'h134 == r_count_50_io_out ? io_r_308_b : _GEN_20487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20489 = 9'h135 == r_count_50_io_out ? io_r_309_b : _GEN_20488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20490 = 9'h136 == r_count_50_io_out ? io_r_310_b : _GEN_20489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20491 = 9'h137 == r_count_50_io_out ? io_r_311_b : _GEN_20490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20492 = 9'h138 == r_count_50_io_out ? io_r_312_b : _GEN_20491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20493 = 9'h139 == r_count_50_io_out ? io_r_313_b : _GEN_20492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20494 = 9'h13a == r_count_50_io_out ? io_r_314_b : _GEN_20493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20495 = 9'h13b == r_count_50_io_out ? io_r_315_b : _GEN_20494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20496 = 9'h13c == r_count_50_io_out ? io_r_316_b : _GEN_20495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20497 = 9'h13d == r_count_50_io_out ? io_r_317_b : _GEN_20496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20498 = 9'h13e == r_count_50_io_out ? io_r_318_b : _GEN_20497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20499 = 9'h13f == r_count_50_io_out ? io_r_319_b : _GEN_20498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20500 = 9'h140 == r_count_50_io_out ? io_r_320_b : _GEN_20499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20501 = 9'h141 == r_count_50_io_out ? io_r_321_b : _GEN_20500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20502 = 9'h142 == r_count_50_io_out ? io_r_322_b : _GEN_20501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20503 = 9'h143 == r_count_50_io_out ? io_r_323_b : _GEN_20502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20504 = 9'h144 == r_count_50_io_out ? io_r_324_b : _GEN_20503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20505 = 9'h145 == r_count_50_io_out ? io_r_325_b : _GEN_20504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20506 = 9'h146 == r_count_50_io_out ? io_r_326_b : _GEN_20505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20507 = 9'h147 == r_count_50_io_out ? io_r_327_b : _GEN_20506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20508 = 9'h148 == r_count_50_io_out ? io_r_328_b : _GEN_20507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20509 = 9'h149 == r_count_50_io_out ? io_r_329_b : _GEN_20508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20510 = 9'h14a == r_count_50_io_out ? io_r_330_b : _GEN_20509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20511 = 9'h14b == r_count_50_io_out ? io_r_331_b : _GEN_20510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20512 = 9'h14c == r_count_50_io_out ? io_r_332_b : _GEN_20511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20513 = 9'h14d == r_count_50_io_out ? io_r_333_b : _GEN_20512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20514 = 9'h14e == r_count_50_io_out ? io_r_334_b : _GEN_20513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20515 = 9'h14f == r_count_50_io_out ? io_r_335_b : _GEN_20514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20516 = 9'h150 == r_count_50_io_out ? io_r_336_b : _GEN_20515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20517 = 9'h151 == r_count_50_io_out ? io_r_337_b : _GEN_20516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20518 = 9'h152 == r_count_50_io_out ? io_r_338_b : _GEN_20517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20519 = 9'h153 == r_count_50_io_out ? io_r_339_b : _GEN_20518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20520 = 9'h154 == r_count_50_io_out ? io_r_340_b : _GEN_20519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20521 = 9'h155 == r_count_50_io_out ? io_r_341_b : _GEN_20520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20522 = 9'h156 == r_count_50_io_out ? io_r_342_b : _GEN_20521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20523 = 9'h157 == r_count_50_io_out ? io_r_343_b : _GEN_20522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20524 = 9'h158 == r_count_50_io_out ? io_r_344_b : _GEN_20523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20525 = 9'h159 == r_count_50_io_out ? io_r_345_b : _GEN_20524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20526 = 9'h15a == r_count_50_io_out ? io_r_346_b : _GEN_20525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20527 = 9'h15b == r_count_50_io_out ? io_r_347_b : _GEN_20526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20528 = 9'h15c == r_count_50_io_out ? io_r_348_b : _GEN_20527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20529 = 9'h15d == r_count_50_io_out ? io_r_349_b : _GEN_20528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20530 = 9'h15e == r_count_50_io_out ? io_r_350_b : _GEN_20529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20531 = 9'h15f == r_count_50_io_out ? io_r_351_b : _GEN_20530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20532 = 9'h160 == r_count_50_io_out ? io_r_352_b : _GEN_20531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20533 = 9'h161 == r_count_50_io_out ? io_r_353_b : _GEN_20532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20534 = 9'h162 == r_count_50_io_out ? io_r_354_b : _GEN_20533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20535 = 9'h163 == r_count_50_io_out ? io_r_355_b : _GEN_20534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20536 = 9'h164 == r_count_50_io_out ? io_r_356_b : _GEN_20535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20537 = 9'h165 == r_count_50_io_out ? io_r_357_b : _GEN_20536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20538 = 9'h166 == r_count_50_io_out ? io_r_358_b : _GEN_20537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20539 = 9'h167 == r_count_50_io_out ? io_r_359_b : _GEN_20538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20540 = 9'h168 == r_count_50_io_out ? io_r_360_b : _GEN_20539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20541 = 9'h169 == r_count_50_io_out ? io_r_361_b : _GEN_20540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20542 = 9'h16a == r_count_50_io_out ? io_r_362_b : _GEN_20541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20543 = 9'h16b == r_count_50_io_out ? io_r_363_b : _GEN_20542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20544 = 9'h16c == r_count_50_io_out ? io_r_364_b : _GEN_20543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20545 = 9'h16d == r_count_50_io_out ? io_r_365_b : _GEN_20544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20546 = 9'h16e == r_count_50_io_out ? io_r_366_b : _GEN_20545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20547 = 9'h16f == r_count_50_io_out ? io_r_367_b : _GEN_20546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20548 = 9'h170 == r_count_50_io_out ? io_r_368_b : _GEN_20547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20549 = 9'h171 == r_count_50_io_out ? io_r_369_b : _GEN_20548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20550 = 9'h172 == r_count_50_io_out ? io_r_370_b : _GEN_20549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20551 = 9'h173 == r_count_50_io_out ? io_r_371_b : _GEN_20550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20552 = 9'h174 == r_count_50_io_out ? io_r_372_b : _GEN_20551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20553 = 9'h175 == r_count_50_io_out ? io_r_373_b : _GEN_20552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20554 = 9'h176 == r_count_50_io_out ? io_r_374_b : _GEN_20553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20555 = 9'h177 == r_count_50_io_out ? io_r_375_b : _GEN_20554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20556 = 9'h178 == r_count_50_io_out ? io_r_376_b : _GEN_20555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20557 = 9'h179 == r_count_50_io_out ? io_r_377_b : _GEN_20556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20558 = 9'h17a == r_count_50_io_out ? io_r_378_b : _GEN_20557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20559 = 9'h17b == r_count_50_io_out ? io_r_379_b : _GEN_20558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20560 = 9'h17c == r_count_50_io_out ? io_r_380_b : _GEN_20559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20561 = 9'h17d == r_count_50_io_out ? io_r_381_b : _GEN_20560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20562 = 9'h17e == r_count_50_io_out ? io_r_382_b : _GEN_20561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20563 = 9'h17f == r_count_50_io_out ? io_r_383_b : _GEN_20562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20564 = 9'h180 == r_count_50_io_out ? io_r_384_b : _GEN_20563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20565 = 9'h181 == r_count_50_io_out ? io_r_385_b : _GEN_20564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20566 = 9'h182 == r_count_50_io_out ? io_r_386_b : _GEN_20565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20567 = 9'h183 == r_count_50_io_out ? io_r_387_b : _GEN_20566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20568 = 9'h184 == r_count_50_io_out ? io_r_388_b : _GEN_20567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20569 = 9'h185 == r_count_50_io_out ? io_r_389_b : _GEN_20568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20570 = 9'h186 == r_count_50_io_out ? io_r_390_b : _GEN_20569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20571 = 9'h187 == r_count_50_io_out ? io_r_391_b : _GEN_20570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20572 = 9'h188 == r_count_50_io_out ? io_r_392_b : _GEN_20571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20573 = 9'h189 == r_count_50_io_out ? io_r_393_b : _GEN_20572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20574 = 9'h18a == r_count_50_io_out ? io_r_394_b : _GEN_20573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20575 = 9'h18b == r_count_50_io_out ? io_r_395_b : _GEN_20574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20576 = 9'h18c == r_count_50_io_out ? io_r_396_b : _GEN_20575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20577 = 9'h18d == r_count_50_io_out ? io_r_397_b : _GEN_20576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20578 = 9'h18e == r_count_50_io_out ? io_r_398_b : _GEN_20577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20581 = 9'h1 == r_count_51_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20582 = 9'h2 == r_count_51_io_out ? io_r_2_b : _GEN_20581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20583 = 9'h3 == r_count_51_io_out ? io_r_3_b : _GEN_20582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20584 = 9'h4 == r_count_51_io_out ? io_r_4_b : _GEN_20583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20585 = 9'h5 == r_count_51_io_out ? io_r_5_b : _GEN_20584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20586 = 9'h6 == r_count_51_io_out ? io_r_6_b : _GEN_20585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20587 = 9'h7 == r_count_51_io_out ? io_r_7_b : _GEN_20586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20588 = 9'h8 == r_count_51_io_out ? io_r_8_b : _GEN_20587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20589 = 9'h9 == r_count_51_io_out ? io_r_9_b : _GEN_20588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20590 = 9'ha == r_count_51_io_out ? io_r_10_b : _GEN_20589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20591 = 9'hb == r_count_51_io_out ? io_r_11_b : _GEN_20590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20592 = 9'hc == r_count_51_io_out ? io_r_12_b : _GEN_20591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20593 = 9'hd == r_count_51_io_out ? io_r_13_b : _GEN_20592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20594 = 9'he == r_count_51_io_out ? io_r_14_b : _GEN_20593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20595 = 9'hf == r_count_51_io_out ? io_r_15_b : _GEN_20594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20596 = 9'h10 == r_count_51_io_out ? io_r_16_b : _GEN_20595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20597 = 9'h11 == r_count_51_io_out ? io_r_17_b : _GEN_20596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20598 = 9'h12 == r_count_51_io_out ? io_r_18_b : _GEN_20597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20599 = 9'h13 == r_count_51_io_out ? io_r_19_b : _GEN_20598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20600 = 9'h14 == r_count_51_io_out ? io_r_20_b : _GEN_20599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20601 = 9'h15 == r_count_51_io_out ? io_r_21_b : _GEN_20600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20602 = 9'h16 == r_count_51_io_out ? io_r_22_b : _GEN_20601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20603 = 9'h17 == r_count_51_io_out ? io_r_23_b : _GEN_20602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20604 = 9'h18 == r_count_51_io_out ? io_r_24_b : _GEN_20603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20605 = 9'h19 == r_count_51_io_out ? io_r_25_b : _GEN_20604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20606 = 9'h1a == r_count_51_io_out ? io_r_26_b : _GEN_20605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20607 = 9'h1b == r_count_51_io_out ? io_r_27_b : _GEN_20606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20608 = 9'h1c == r_count_51_io_out ? io_r_28_b : _GEN_20607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20609 = 9'h1d == r_count_51_io_out ? io_r_29_b : _GEN_20608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20610 = 9'h1e == r_count_51_io_out ? io_r_30_b : _GEN_20609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20611 = 9'h1f == r_count_51_io_out ? io_r_31_b : _GEN_20610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20612 = 9'h20 == r_count_51_io_out ? io_r_32_b : _GEN_20611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20613 = 9'h21 == r_count_51_io_out ? io_r_33_b : _GEN_20612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20614 = 9'h22 == r_count_51_io_out ? io_r_34_b : _GEN_20613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20615 = 9'h23 == r_count_51_io_out ? io_r_35_b : _GEN_20614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20616 = 9'h24 == r_count_51_io_out ? io_r_36_b : _GEN_20615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20617 = 9'h25 == r_count_51_io_out ? io_r_37_b : _GEN_20616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20618 = 9'h26 == r_count_51_io_out ? io_r_38_b : _GEN_20617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20619 = 9'h27 == r_count_51_io_out ? io_r_39_b : _GEN_20618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20620 = 9'h28 == r_count_51_io_out ? io_r_40_b : _GEN_20619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20621 = 9'h29 == r_count_51_io_out ? io_r_41_b : _GEN_20620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20622 = 9'h2a == r_count_51_io_out ? io_r_42_b : _GEN_20621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20623 = 9'h2b == r_count_51_io_out ? io_r_43_b : _GEN_20622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20624 = 9'h2c == r_count_51_io_out ? io_r_44_b : _GEN_20623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20625 = 9'h2d == r_count_51_io_out ? io_r_45_b : _GEN_20624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20626 = 9'h2e == r_count_51_io_out ? io_r_46_b : _GEN_20625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20627 = 9'h2f == r_count_51_io_out ? io_r_47_b : _GEN_20626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20628 = 9'h30 == r_count_51_io_out ? io_r_48_b : _GEN_20627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20629 = 9'h31 == r_count_51_io_out ? io_r_49_b : _GEN_20628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20630 = 9'h32 == r_count_51_io_out ? io_r_50_b : _GEN_20629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20631 = 9'h33 == r_count_51_io_out ? io_r_51_b : _GEN_20630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20632 = 9'h34 == r_count_51_io_out ? io_r_52_b : _GEN_20631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20633 = 9'h35 == r_count_51_io_out ? io_r_53_b : _GEN_20632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20634 = 9'h36 == r_count_51_io_out ? io_r_54_b : _GEN_20633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20635 = 9'h37 == r_count_51_io_out ? io_r_55_b : _GEN_20634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20636 = 9'h38 == r_count_51_io_out ? io_r_56_b : _GEN_20635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20637 = 9'h39 == r_count_51_io_out ? io_r_57_b : _GEN_20636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20638 = 9'h3a == r_count_51_io_out ? io_r_58_b : _GEN_20637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20639 = 9'h3b == r_count_51_io_out ? io_r_59_b : _GEN_20638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20640 = 9'h3c == r_count_51_io_out ? io_r_60_b : _GEN_20639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20641 = 9'h3d == r_count_51_io_out ? io_r_61_b : _GEN_20640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20642 = 9'h3e == r_count_51_io_out ? io_r_62_b : _GEN_20641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20643 = 9'h3f == r_count_51_io_out ? io_r_63_b : _GEN_20642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20644 = 9'h40 == r_count_51_io_out ? io_r_64_b : _GEN_20643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20645 = 9'h41 == r_count_51_io_out ? io_r_65_b : _GEN_20644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20646 = 9'h42 == r_count_51_io_out ? io_r_66_b : _GEN_20645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20647 = 9'h43 == r_count_51_io_out ? io_r_67_b : _GEN_20646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20648 = 9'h44 == r_count_51_io_out ? io_r_68_b : _GEN_20647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20649 = 9'h45 == r_count_51_io_out ? io_r_69_b : _GEN_20648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20650 = 9'h46 == r_count_51_io_out ? io_r_70_b : _GEN_20649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20651 = 9'h47 == r_count_51_io_out ? io_r_71_b : _GEN_20650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20652 = 9'h48 == r_count_51_io_out ? io_r_72_b : _GEN_20651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20653 = 9'h49 == r_count_51_io_out ? io_r_73_b : _GEN_20652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20654 = 9'h4a == r_count_51_io_out ? io_r_74_b : _GEN_20653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20655 = 9'h4b == r_count_51_io_out ? io_r_75_b : _GEN_20654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20656 = 9'h4c == r_count_51_io_out ? io_r_76_b : _GEN_20655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20657 = 9'h4d == r_count_51_io_out ? io_r_77_b : _GEN_20656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20658 = 9'h4e == r_count_51_io_out ? io_r_78_b : _GEN_20657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20659 = 9'h4f == r_count_51_io_out ? io_r_79_b : _GEN_20658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20660 = 9'h50 == r_count_51_io_out ? io_r_80_b : _GEN_20659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20661 = 9'h51 == r_count_51_io_out ? io_r_81_b : _GEN_20660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20662 = 9'h52 == r_count_51_io_out ? io_r_82_b : _GEN_20661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20663 = 9'h53 == r_count_51_io_out ? io_r_83_b : _GEN_20662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20664 = 9'h54 == r_count_51_io_out ? io_r_84_b : _GEN_20663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20665 = 9'h55 == r_count_51_io_out ? io_r_85_b : _GEN_20664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20666 = 9'h56 == r_count_51_io_out ? io_r_86_b : _GEN_20665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20667 = 9'h57 == r_count_51_io_out ? io_r_87_b : _GEN_20666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20668 = 9'h58 == r_count_51_io_out ? io_r_88_b : _GEN_20667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20669 = 9'h59 == r_count_51_io_out ? io_r_89_b : _GEN_20668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20670 = 9'h5a == r_count_51_io_out ? io_r_90_b : _GEN_20669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20671 = 9'h5b == r_count_51_io_out ? io_r_91_b : _GEN_20670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20672 = 9'h5c == r_count_51_io_out ? io_r_92_b : _GEN_20671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20673 = 9'h5d == r_count_51_io_out ? io_r_93_b : _GEN_20672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20674 = 9'h5e == r_count_51_io_out ? io_r_94_b : _GEN_20673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20675 = 9'h5f == r_count_51_io_out ? io_r_95_b : _GEN_20674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20676 = 9'h60 == r_count_51_io_out ? io_r_96_b : _GEN_20675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20677 = 9'h61 == r_count_51_io_out ? io_r_97_b : _GEN_20676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20678 = 9'h62 == r_count_51_io_out ? io_r_98_b : _GEN_20677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20679 = 9'h63 == r_count_51_io_out ? io_r_99_b : _GEN_20678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20680 = 9'h64 == r_count_51_io_out ? io_r_100_b : _GEN_20679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20681 = 9'h65 == r_count_51_io_out ? io_r_101_b : _GEN_20680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20682 = 9'h66 == r_count_51_io_out ? io_r_102_b : _GEN_20681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20683 = 9'h67 == r_count_51_io_out ? io_r_103_b : _GEN_20682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20684 = 9'h68 == r_count_51_io_out ? io_r_104_b : _GEN_20683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20685 = 9'h69 == r_count_51_io_out ? io_r_105_b : _GEN_20684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20686 = 9'h6a == r_count_51_io_out ? io_r_106_b : _GEN_20685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20687 = 9'h6b == r_count_51_io_out ? io_r_107_b : _GEN_20686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20688 = 9'h6c == r_count_51_io_out ? io_r_108_b : _GEN_20687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20689 = 9'h6d == r_count_51_io_out ? io_r_109_b : _GEN_20688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20690 = 9'h6e == r_count_51_io_out ? io_r_110_b : _GEN_20689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20691 = 9'h6f == r_count_51_io_out ? io_r_111_b : _GEN_20690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20692 = 9'h70 == r_count_51_io_out ? io_r_112_b : _GEN_20691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20693 = 9'h71 == r_count_51_io_out ? io_r_113_b : _GEN_20692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20694 = 9'h72 == r_count_51_io_out ? io_r_114_b : _GEN_20693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20695 = 9'h73 == r_count_51_io_out ? io_r_115_b : _GEN_20694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20696 = 9'h74 == r_count_51_io_out ? io_r_116_b : _GEN_20695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20697 = 9'h75 == r_count_51_io_out ? io_r_117_b : _GEN_20696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20698 = 9'h76 == r_count_51_io_out ? io_r_118_b : _GEN_20697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20699 = 9'h77 == r_count_51_io_out ? io_r_119_b : _GEN_20698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20700 = 9'h78 == r_count_51_io_out ? io_r_120_b : _GEN_20699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20701 = 9'h79 == r_count_51_io_out ? io_r_121_b : _GEN_20700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20702 = 9'h7a == r_count_51_io_out ? io_r_122_b : _GEN_20701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20703 = 9'h7b == r_count_51_io_out ? io_r_123_b : _GEN_20702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20704 = 9'h7c == r_count_51_io_out ? io_r_124_b : _GEN_20703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20705 = 9'h7d == r_count_51_io_out ? io_r_125_b : _GEN_20704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20706 = 9'h7e == r_count_51_io_out ? io_r_126_b : _GEN_20705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20707 = 9'h7f == r_count_51_io_out ? io_r_127_b : _GEN_20706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20708 = 9'h80 == r_count_51_io_out ? io_r_128_b : _GEN_20707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20709 = 9'h81 == r_count_51_io_out ? io_r_129_b : _GEN_20708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20710 = 9'h82 == r_count_51_io_out ? io_r_130_b : _GEN_20709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20711 = 9'h83 == r_count_51_io_out ? io_r_131_b : _GEN_20710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20712 = 9'h84 == r_count_51_io_out ? io_r_132_b : _GEN_20711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20713 = 9'h85 == r_count_51_io_out ? io_r_133_b : _GEN_20712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20714 = 9'h86 == r_count_51_io_out ? io_r_134_b : _GEN_20713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20715 = 9'h87 == r_count_51_io_out ? io_r_135_b : _GEN_20714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20716 = 9'h88 == r_count_51_io_out ? io_r_136_b : _GEN_20715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20717 = 9'h89 == r_count_51_io_out ? io_r_137_b : _GEN_20716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20718 = 9'h8a == r_count_51_io_out ? io_r_138_b : _GEN_20717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20719 = 9'h8b == r_count_51_io_out ? io_r_139_b : _GEN_20718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20720 = 9'h8c == r_count_51_io_out ? io_r_140_b : _GEN_20719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20721 = 9'h8d == r_count_51_io_out ? io_r_141_b : _GEN_20720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20722 = 9'h8e == r_count_51_io_out ? io_r_142_b : _GEN_20721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20723 = 9'h8f == r_count_51_io_out ? io_r_143_b : _GEN_20722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20724 = 9'h90 == r_count_51_io_out ? io_r_144_b : _GEN_20723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20725 = 9'h91 == r_count_51_io_out ? io_r_145_b : _GEN_20724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20726 = 9'h92 == r_count_51_io_out ? io_r_146_b : _GEN_20725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20727 = 9'h93 == r_count_51_io_out ? io_r_147_b : _GEN_20726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20728 = 9'h94 == r_count_51_io_out ? io_r_148_b : _GEN_20727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20729 = 9'h95 == r_count_51_io_out ? io_r_149_b : _GEN_20728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20730 = 9'h96 == r_count_51_io_out ? io_r_150_b : _GEN_20729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20731 = 9'h97 == r_count_51_io_out ? io_r_151_b : _GEN_20730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20732 = 9'h98 == r_count_51_io_out ? io_r_152_b : _GEN_20731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20733 = 9'h99 == r_count_51_io_out ? io_r_153_b : _GEN_20732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20734 = 9'h9a == r_count_51_io_out ? io_r_154_b : _GEN_20733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20735 = 9'h9b == r_count_51_io_out ? io_r_155_b : _GEN_20734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20736 = 9'h9c == r_count_51_io_out ? io_r_156_b : _GEN_20735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20737 = 9'h9d == r_count_51_io_out ? io_r_157_b : _GEN_20736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20738 = 9'h9e == r_count_51_io_out ? io_r_158_b : _GEN_20737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20739 = 9'h9f == r_count_51_io_out ? io_r_159_b : _GEN_20738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20740 = 9'ha0 == r_count_51_io_out ? io_r_160_b : _GEN_20739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20741 = 9'ha1 == r_count_51_io_out ? io_r_161_b : _GEN_20740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20742 = 9'ha2 == r_count_51_io_out ? io_r_162_b : _GEN_20741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20743 = 9'ha3 == r_count_51_io_out ? io_r_163_b : _GEN_20742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20744 = 9'ha4 == r_count_51_io_out ? io_r_164_b : _GEN_20743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20745 = 9'ha5 == r_count_51_io_out ? io_r_165_b : _GEN_20744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20746 = 9'ha6 == r_count_51_io_out ? io_r_166_b : _GEN_20745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20747 = 9'ha7 == r_count_51_io_out ? io_r_167_b : _GEN_20746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20748 = 9'ha8 == r_count_51_io_out ? io_r_168_b : _GEN_20747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20749 = 9'ha9 == r_count_51_io_out ? io_r_169_b : _GEN_20748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20750 = 9'haa == r_count_51_io_out ? io_r_170_b : _GEN_20749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20751 = 9'hab == r_count_51_io_out ? io_r_171_b : _GEN_20750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20752 = 9'hac == r_count_51_io_out ? io_r_172_b : _GEN_20751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20753 = 9'had == r_count_51_io_out ? io_r_173_b : _GEN_20752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20754 = 9'hae == r_count_51_io_out ? io_r_174_b : _GEN_20753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20755 = 9'haf == r_count_51_io_out ? io_r_175_b : _GEN_20754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20756 = 9'hb0 == r_count_51_io_out ? io_r_176_b : _GEN_20755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20757 = 9'hb1 == r_count_51_io_out ? io_r_177_b : _GEN_20756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20758 = 9'hb2 == r_count_51_io_out ? io_r_178_b : _GEN_20757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20759 = 9'hb3 == r_count_51_io_out ? io_r_179_b : _GEN_20758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20760 = 9'hb4 == r_count_51_io_out ? io_r_180_b : _GEN_20759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20761 = 9'hb5 == r_count_51_io_out ? io_r_181_b : _GEN_20760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20762 = 9'hb6 == r_count_51_io_out ? io_r_182_b : _GEN_20761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20763 = 9'hb7 == r_count_51_io_out ? io_r_183_b : _GEN_20762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20764 = 9'hb8 == r_count_51_io_out ? io_r_184_b : _GEN_20763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20765 = 9'hb9 == r_count_51_io_out ? io_r_185_b : _GEN_20764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20766 = 9'hba == r_count_51_io_out ? io_r_186_b : _GEN_20765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20767 = 9'hbb == r_count_51_io_out ? io_r_187_b : _GEN_20766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20768 = 9'hbc == r_count_51_io_out ? io_r_188_b : _GEN_20767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20769 = 9'hbd == r_count_51_io_out ? io_r_189_b : _GEN_20768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20770 = 9'hbe == r_count_51_io_out ? io_r_190_b : _GEN_20769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20771 = 9'hbf == r_count_51_io_out ? io_r_191_b : _GEN_20770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20772 = 9'hc0 == r_count_51_io_out ? io_r_192_b : _GEN_20771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20773 = 9'hc1 == r_count_51_io_out ? io_r_193_b : _GEN_20772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20774 = 9'hc2 == r_count_51_io_out ? io_r_194_b : _GEN_20773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20775 = 9'hc3 == r_count_51_io_out ? io_r_195_b : _GEN_20774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20776 = 9'hc4 == r_count_51_io_out ? io_r_196_b : _GEN_20775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20777 = 9'hc5 == r_count_51_io_out ? io_r_197_b : _GEN_20776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20778 = 9'hc6 == r_count_51_io_out ? io_r_198_b : _GEN_20777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20779 = 9'hc7 == r_count_51_io_out ? io_r_199_b : _GEN_20778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20780 = 9'hc8 == r_count_51_io_out ? io_r_200_b : _GEN_20779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20781 = 9'hc9 == r_count_51_io_out ? io_r_201_b : _GEN_20780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20782 = 9'hca == r_count_51_io_out ? io_r_202_b : _GEN_20781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20783 = 9'hcb == r_count_51_io_out ? io_r_203_b : _GEN_20782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20784 = 9'hcc == r_count_51_io_out ? io_r_204_b : _GEN_20783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20785 = 9'hcd == r_count_51_io_out ? io_r_205_b : _GEN_20784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20786 = 9'hce == r_count_51_io_out ? io_r_206_b : _GEN_20785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20787 = 9'hcf == r_count_51_io_out ? io_r_207_b : _GEN_20786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20788 = 9'hd0 == r_count_51_io_out ? io_r_208_b : _GEN_20787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20789 = 9'hd1 == r_count_51_io_out ? io_r_209_b : _GEN_20788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20790 = 9'hd2 == r_count_51_io_out ? io_r_210_b : _GEN_20789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20791 = 9'hd3 == r_count_51_io_out ? io_r_211_b : _GEN_20790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20792 = 9'hd4 == r_count_51_io_out ? io_r_212_b : _GEN_20791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20793 = 9'hd5 == r_count_51_io_out ? io_r_213_b : _GEN_20792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20794 = 9'hd6 == r_count_51_io_out ? io_r_214_b : _GEN_20793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20795 = 9'hd7 == r_count_51_io_out ? io_r_215_b : _GEN_20794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20796 = 9'hd8 == r_count_51_io_out ? io_r_216_b : _GEN_20795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20797 = 9'hd9 == r_count_51_io_out ? io_r_217_b : _GEN_20796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20798 = 9'hda == r_count_51_io_out ? io_r_218_b : _GEN_20797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20799 = 9'hdb == r_count_51_io_out ? io_r_219_b : _GEN_20798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20800 = 9'hdc == r_count_51_io_out ? io_r_220_b : _GEN_20799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20801 = 9'hdd == r_count_51_io_out ? io_r_221_b : _GEN_20800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20802 = 9'hde == r_count_51_io_out ? io_r_222_b : _GEN_20801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20803 = 9'hdf == r_count_51_io_out ? io_r_223_b : _GEN_20802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20804 = 9'he0 == r_count_51_io_out ? io_r_224_b : _GEN_20803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20805 = 9'he1 == r_count_51_io_out ? io_r_225_b : _GEN_20804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20806 = 9'he2 == r_count_51_io_out ? io_r_226_b : _GEN_20805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20807 = 9'he3 == r_count_51_io_out ? io_r_227_b : _GEN_20806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20808 = 9'he4 == r_count_51_io_out ? io_r_228_b : _GEN_20807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20809 = 9'he5 == r_count_51_io_out ? io_r_229_b : _GEN_20808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20810 = 9'he6 == r_count_51_io_out ? io_r_230_b : _GEN_20809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20811 = 9'he7 == r_count_51_io_out ? io_r_231_b : _GEN_20810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20812 = 9'he8 == r_count_51_io_out ? io_r_232_b : _GEN_20811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20813 = 9'he9 == r_count_51_io_out ? io_r_233_b : _GEN_20812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20814 = 9'hea == r_count_51_io_out ? io_r_234_b : _GEN_20813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20815 = 9'heb == r_count_51_io_out ? io_r_235_b : _GEN_20814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20816 = 9'hec == r_count_51_io_out ? io_r_236_b : _GEN_20815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20817 = 9'hed == r_count_51_io_out ? io_r_237_b : _GEN_20816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20818 = 9'hee == r_count_51_io_out ? io_r_238_b : _GEN_20817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20819 = 9'hef == r_count_51_io_out ? io_r_239_b : _GEN_20818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20820 = 9'hf0 == r_count_51_io_out ? io_r_240_b : _GEN_20819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20821 = 9'hf1 == r_count_51_io_out ? io_r_241_b : _GEN_20820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20822 = 9'hf2 == r_count_51_io_out ? io_r_242_b : _GEN_20821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20823 = 9'hf3 == r_count_51_io_out ? io_r_243_b : _GEN_20822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20824 = 9'hf4 == r_count_51_io_out ? io_r_244_b : _GEN_20823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20825 = 9'hf5 == r_count_51_io_out ? io_r_245_b : _GEN_20824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20826 = 9'hf6 == r_count_51_io_out ? io_r_246_b : _GEN_20825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20827 = 9'hf7 == r_count_51_io_out ? io_r_247_b : _GEN_20826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20828 = 9'hf8 == r_count_51_io_out ? io_r_248_b : _GEN_20827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20829 = 9'hf9 == r_count_51_io_out ? io_r_249_b : _GEN_20828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20830 = 9'hfa == r_count_51_io_out ? io_r_250_b : _GEN_20829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20831 = 9'hfb == r_count_51_io_out ? io_r_251_b : _GEN_20830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20832 = 9'hfc == r_count_51_io_out ? io_r_252_b : _GEN_20831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20833 = 9'hfd == r_count_51_io_out ? io_r_253_b : _GEN_20832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20834 = 9'hfe == r_count_51_io_out ? io_r_254_b : _GEN_20833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20835 = 9'hff == r_count_51_io_out ? io_r_255_b : _GEN_20834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20836 = 9'h100 == r_count_51_io_out ? io_r_256_b : _GEN_20835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20837 = 9'h101 == r_count_51_io_out ? io_r_257_b : _GEN_20836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20838 = 9'h102 == r_count_51_io_out ? io_r_258_b : _GEN_20837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20839 = 9'h103 == r_count_51_io_out ? io_r_259_b : _GEN_20838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20840 = 9'h104 == r_count_51_io_out ? io_r_260_b : _GEN_20839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20841 = 9'h105 == r_count_51_io_out ? io_r_261_b : _GEN_20840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20842 = 9'h106 == r_count_51_io_out ? io_r_262_b : _GEN_20841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20843 = 9'h107 == r_count_51_io_out ? io_r_263_b : _GEN_20842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20844 = 9'h108 == r_count_51_io_out ? io_r_264_b : _GEN_20843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20845 = 9'h109 == r_count_51_io_out ? io_r_265_b : _GEN_20844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20846 = 9'h10a == r_count_51_io_out ? io_r_266_b : _GEN_20845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20847 = 9'h10b == r_count_51_io_out ? io_r_267_b : _GEN_20846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20848 = 9'h10c == r_count_51_io_out ? io_r_268_b : _GEN_20847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20849 = 9'h10d == r_count_51_io_out ? io_r_269_b : _GEN_20848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20850 = 9'h10e == r_count_51_io_out ? io_r_270_b : _GEN_20849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20851 = 9'h10f == r_count_51_io_out ? io_r_271_b : _GEN_20850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20852 = 9'h110 == r_count_51_io_out ? io_r_272_b : _GEN_20851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20853 = 9'h111 == r_count_51_io_out ? io_r_273_b : _GEN_20852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20854 = 9'h112 == r_count_51_io_out ? io_r_274_b : _GEN_20853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20855 = 9'h113 == r_count_51_io_out ? io_r_275_b : _GEN_20854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20856 = 9'h114 == r_count_51_io_out ? io_r_276_b : _GEN_20855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20857 = 9'h115 == r_count_51_io_out ? io_r_277_b : _GEN_20856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20858 = 9'h116 == r_count_51_io_out ? io_r_278_b : _GEN_20857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20859 = 9'h117 == r_count_51_io_out ? io_r_279_b : _GEN_20858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20860 = 9'h118 == r_count_51_io_out ? io_r_280_b : _GEN_20859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20861 = 9'h119 == r_count_51_io_out ? io_r_281_b : _GEN_20860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20862 = 9'h11a == r_count_51_io_out ? io_r_282_b : _GEN_20861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20863 = 9'h11b == r_count_51_io_out ? io_r_283_b : _GEN_20862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20864 = 9'h11c == r_count_51_io_out ? io_r_284_b : _GEN_20863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20865 = 9'h11d == r_count_51_io_out ? io_r_285_b : _GEN_20864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20866 = 9'h11e == r_count_51_io_out ? io_r_286_b : _GEN_20865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20867 = 9'h11f == r_count_51_io_out ? io_r_287_b : _GEN_20866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20868 = 9'h120 == r_count_51_io_out ? io_r_288_b : _GEN_20867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20869 = 9'h121 == r_count_51_io_out ? io_r_289_b : _GEN_20868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20870 = 9'h122 == r_count_51_io_out ? io_r_290_b : _GEN_20869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20871 = 9'h123 == r_count_51_io_out ? io_r_291_b : _GEN_20870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20872 = 9'h124 == r_count_51_io_out ? io_r_292_b : _GEN_20871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20873 = 9'h125 == r_count_51_io_out ? io_r_293_b : _GEN_20872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20874 = 9'h126 == r_count_51_io_out ? io_r_294_b : _GEN_20873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20875 = 9'h127 == r_count_51_io_out ? io_r_295_b : _GEN_20874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20876 = 9'h128 == r_count_51_io_out ? io_r_296_b : _GEN_20875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20877 = 9'h129 == r_count_51_io_out ? io_r_297_b : _GEN_20876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20878 = 9'h12a == r_count_51_io_out ? io_r_298_b : _GEN_20877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20879 = 9'h12b == r_count_51_io_out ? io_r_299_b : _GEN_20878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20880 = 9'h12c == r_count_51_io_out ? io_r_300_b : _GEN_20879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20881 = 9'h12d == r_count_51_io_out ? io_r_301_b : _GEN_20880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20882 = 9'h12e == r_count_51_io_out ? io_r_302_b : _GEN_20881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20883 = 9'h12f == r_count_51_io_out ? io_r_303_b : _GEN_20882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20884 = 9'h130 == r_count_51_io_out ? io_r_304_b : _GEN_20883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20885 = 9'h131 == r_count_51_io_out ? io_r_305_b : _GEN_20884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20886 = 9'h132 == r_count_51_io_out ? io_r_306_b : _GEN_20885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20887 = 9'h133 == r_count_51_io_out ? io_r_307_b : _GEN_20886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20888 = 9'h134 == r_count_51_io_out ? io_r_308_b : _GEN_20887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20889 = 9'h135 == r_count_51_io_out ? io_r_309_b : _GEN_20888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20890 = 9'h136 == r_count_51_io_out ? io_r_310_b : _GEN_20889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20891 = 9'h137 == r_count_51_io_out ? io_r_311_b : _GEN_20890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20892 = 9'h138 == r_count_51_io_out ? io_r_312_b : _GEN_20891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20893 = 9'h139 == r_count_51_io_out ? io_r_313_b : _GEN_20892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20894 = 9'h13a == r_count_51_io_out ? io_r_314_b : _GEN_20893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20895 = 9'h13b == r_count_51_io_out ? io_r_315_b : _GEN_20894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20896 = 9'h13c == r_count_51_io_out ? io_r_316_b : _GEN_20895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20897 = 9'h13d == r_count_51_io_out ? io_r_317_b : _GEN_20896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20898 = 9'h13e == r_count_51_io_out ? io_r_318_b : _GEN_20897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20899 = 9'h13f == r_count_51_io_out ? io_r_319_b : _GEN_20898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20900 = 9'h140 == r_count_51_io_out ? io_r_320_b : _GEN_20899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20901 = 9'h141 == r_count_51_io_out ? io_r_321_b : _GEN_20900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20902 = 9'h142 == r_count_51_io_out ? io_r_322_b : _GEN_20901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20903 = 9'h143 == r_count_51_io_out ? io_r_323_b : _GEN_20902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20904 = 9'h144 == r_count_51_io_out ? io_r_324_b : _GEN_20903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20905 = 9'h145 == r_count_51_io_out ? io_r_325_b : _GEN_20904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20906 = 9'h146 == r_count_51_io_out ? io_r_326_b : _GEN_20905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20907 = 9'h147 == r_count_51_io_out ? io_r_327_b : _GEN_20906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20908 = 9'h148 == r_count_51_io_out ? io_r_328_b : _GEN_20907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20909 = 9'h149 == r_count_51_io_out ? io_r_329_b : _GEN_20908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20910 = 9'h14a == r_count_51_io_out ? io_r_330_b : _GEN_20909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20911 = 9'h14b == r_count_51_io_out ? io_r_331_b : _GEN_20910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20912 = 9'h14c == r_count_51_io_out ? io_r_332_b : _GEN_20911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20913 = 9'h14d == r_count_51_io_out ? io_r_333_b : _GEN_20912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20914 = 9'h14e == r_count_51_io_out ? io_r_334_b : _GEN_20913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20915 = 9'h14f == r_count_51_io_out ? io_r_335_b : _GEN_20914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20916 = 9'h150 == r_count_51_io_out ? io_r_336_b : _GEN_20915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20917 = 9'h151 == r_count_51_io_out ? io_r_337_b : _GEN_20916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20918 = 9'h152 == r_count_51_io_out ? io_r_338_b : _GEN_20917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20919 = 9'h153 == r_count_51_io_out ? io_r_339_b : _GEN_20918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20920 = 9'h154 == r_count_51_io_out ? io_r_340_b : _GEN_20919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20921 = 9'h155 == r_count_51_io_out ? io_r_341_b : _GEN_20920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20922 = 9'h156 == r_count_51_io_out ? io_r_342_b : _GEN_20921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20923 = 9'h157 == r_count_51_io_out ? io_r_343_b : _GEN_20922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20924 = 9'h158 == r_count_51_io_out ? io_r_344_b : _GEN_20923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20925 = 9'h159 == r_count_51_io_out ? io_r_345_b : _GEN_20924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20926 = 9'h15a == r_count_51_io_out ? io_r_346_b : _GEN_20925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20927 = 9'h15b == r_count_51_io_out ? io_r_347_b : _GEN_20926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20928 = 9'h15c == r_count_51_io_out ? io_r_348_b : _GEN_20927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20929 = 9'h15d == r_count_51_io_out ? io_r_349_b : _GEN_20928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20930 = 9'h15e == r_count_51_io_out ? io_r_350_b : _GEN_20929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20931 = 9'h15f == r_count_51_io_out ? io_r_351_b : _GEN_20930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20932 = 9'h160 == r_count_51_io_out ? io_r_352_b : _GEN_20931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20933 = 9'h161 == r_count_51_io_out ? io_r_353_b : _GEN_20932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20934 = 9'h162 == r_count_51_io_out ? io_r_354_b : _GEN_20933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20935 = 9'h163 == r_count_51_io_out ? io_r_355_b : _GEN_20934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20936 = 9'h164 == r_count_51_io_out ? io_r_356_b : _GEN_20935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20937 = 9'h165 == r_count_51_io_out ? io_r_357_b : _GEN_20936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20938 = 9'h166 == r_count_51_io_out ? io_r_358_b : _GEN_20937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20939 = 9'h167 == r_count_51_io_out ? io_r_359_b : _GEN_20938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20940 = 9'h168 == r_count_51_io_out ? io_r_360_b : _GEN_20939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20941 = 9'h169 == r_count_51_io_out ? io_r_361_b : _GEN_20940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20942 = 9'h16a == r_count_51_io_out ? io_r_362_b : _GEN_20941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20943 = 9'h16b == r_count_51_io_out ? io_r_363_b : _GEN_20942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20944 = 9'h16c == r_count_51_io_out ? io_r_364_b : _GEN_20943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20945 = 9'h16d == r_count_51_io_out ? io_r_365_b : _GEN_20944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20946 = 9'h16e == r_count_51_io_out ? io_r_366_b : _GEN_20945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20947 = 9'h16f == r_count_51_io_out ? io_r_367_b : _GEN_20946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20948 = 9'h170 == r_count_51_io_out ? io_r_368_b : _GEN_20947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20949 = 9'h171 == r_count_51_io_out ? io_r_369_b : _GEN_20948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20950 = 9'h172 == r_count_51_io_out ? io_r_370_b : _GEN_20949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20951 = 9'h173 == r_count_51_io_out ? io_r_371_b : _GEN_20950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20952 = 9'h174 == r_count_51_io_out ? io_r_372_b : _GEN_20951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20953 = 9'h175 == r_count_51_io_out ? io_r_373_b : _GEN_20952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20954 = 9'h176 == r_count_51_io_out ? io_r_374_b : _GEN_20953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20955 = 9'h177 == r_count_51_io_out ? io_r_375_b : _GEN_20954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20956 = 9'h178 == r_count_51_io_out ? io_r_376_b : _GEN_20955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20957 = 9'h179 == r_count_51_io_out ? io_r_377_b : _GEN_20956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20958 = 9'h17a == r_count_51_io_out ? io_r_378_b : _GEN_20957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20959 = 9'h17b == r_count_51_io_out ? io_r_379_b : _GEN_20958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20960 = 9'h17c == r_count_51_io_out ? io_r_380_b : _GEN_20959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20961 = 9'h17d == r_count_51_io_out ? io_r_381_b : _GEN_20960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20962 = 9'h17e == r_count_51_io_out ? io_r_382_b : _GEN_20961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20963 = 9'h17f == r_count_51_io_out ? io_r_383_b : _GEN_20962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20964 = 9'h180 == r_count_51_io_out ? io_r_384_b : _GEN_20963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20965 = 9'h181 == r_count_51_io_out ? io_r_385_b : _GEN_20964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20966 = 9'h182 == r_count_51_io_out ? io_r_386_b : _GEN_20965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20967 = 9'h183 == r_count_51_io_out ? io_r_387_b : _GEN_20966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20968 = 9'h184 == r_count_51_io_out ? io_r_388_b : _GEN_20967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20969 = 9'h185 == r_count_51_io_out ? io_r_389_b : _GEN_20968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20970 = 9'h186 == r_count_51_io_out ? io_r_390_b : _GEN_20969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20971 = 9'h187 == r_count_51_io_out ? io_r_391_b : _GEN_20970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20972 = 9'h188 == r_count_51_io_out ? io_r_392_b : _GEN_20971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20973 = 9'h189 == r_count_51_io_out ? io_r_393_b : _GEN_20972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20974 = 9'h18a == r_count_51_io_out ? io_r_394_b : _GEN_20973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20975 = 9'h18b == r_count_51_io_out ? io_r_395_b : _GEN_20974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20976 = 9'h18c == r_count_51_io_out ? io_r_396_b : _GEN_20975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20977 = 9'h18d == r_count_51_io_out ? io_r_397_b : _GEN_20976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20978 = 9'h18e == r_count_51_io_out ? io_r_398_b : _GEN_20977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20981 = 9'h1 == r_count_52_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20982 = 9'h2 == r_count_52_io_out ? io_r_2_b : _GEN_20981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20983 = 9'h3 == r_count_52_io_out ? io_r_3_b : _GEN_20982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20984 = 9'h4 == r_count_52_io_out ? io_r_4_b : _GEN_20983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20985 = 9'h5 == r_count_52_io_out ? io_r_5_b : _GEN_20984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20986 = 9'h6 == r_count_52_io_out ? io_r_6_b : _GEN_20985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20987 = 9'h7 == r_count_52_io_out ? io_r_7_b : _GEN_20986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20988 = 9'h8 == r_count_52_io_out ? io_r_8_b : _GEN_20987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20989 = 9'h9 == r_count_52_io_out ? io_r_9_b : _GEN_20988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20990 = 9'ha == r_count_52_io_out ? io_r_10_b : _GEN_20989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20991 = 9'hb == r_count_52_io_out ? io_r_11_b : _GEN_20990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20992 = 9'hc == r_count_52_io_out ? io_r_12_b : _GEN_20991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20993 = 9'hd == r_count_52_io_out ? io_r_13_b : _GEN_20992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20994 = 9'he == r_count_52_io_out ? io_r_14_b : _GEN_20993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20995 = 9'hf == r_count_52_io_out ? io_r_15_b : _GEN_20994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20996 = 9'h10 == r_count_52_io_out ? io_r_16_b : _GEN_20995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20997 = 9'h11 == r_count_52_io_out ? io_r_17_b : _GEN_20996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20998 = 9'h12 == r_count_52_io_out ? io_r_18_b : _GEN_20997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20999 = 9'h13 == r_count_52_io_out ? io_r_19_b : _GEN_20998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21000 = 9'h14 == r_count_52_io_out ? io_r_20_b : _GEN_20999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21001 = 9'h15 == r_count_52_io_out ? io_r_21_b : _GEN_21000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21002 = 9'h16 == r_count_52_io_out ? io_r_22_b : _GEN_21001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21003 = 9'h17 == r_count_52_io_out ? io_r_23_b : _GEN_21002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21004 = 9'h18 == r_count_52_io_out ? io_r_24_b : _GEN_21003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21005 = 9'h19 == r_count_52_io_out ? io_r_25_b : _GEN_21004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21006 = 9'h1a == r_count_52_io_out ? io_r_26_b : _GEN_21005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21007 = 9'h1b == r_count_52_io_out ? io_r_27_b : _GEN_21006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21008 = 9'h1c == r_count_52_io_out ? io_r_28_b : _GEN_21007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21009 = 9'h1d == r_count_52_io_out ? io_r_29_b : _GEN_21008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21010 = 9'h1e == r_count_52_io_out ? io_r_30_b : _GEN_21009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21011 = 9'h1f == r_count_52_io_out ? io_r_31_b : _GEN_21010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21012 = 9'h20 == r_count_52_io_out ? io_r_32_b : _GEN_21011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21013 = 9'h21 == r_count_52_io_out ? io_r_33_b : _GEN_21012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21014 = 9'h22 == r_count_52_io_out ? io_r_34_b : _GEN_21013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21015 = 9'h23 == r_count_52_io_out ? io_r_35_b : _GEN_21014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21016 = 9'h24 == r_count_52_io_out ? io_r_36_b : _GEN_21015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21017 = 9'h25 == r_count_52_io_out ? io_r_37_b : _GEN_21016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21018 = 9'h26 == r_count_52_io_out ? io_r_38_b : _GEN_21017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21019 = 9'h27 == r_count_52_io_out ? io_r_39_b : _GEN_21018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21020 = 9'h28 == r_count_52_io_out ? io_r_40_b : _GEN_21019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21021 = 9'h29 == r_count_52_io_out ? io_r_41_b : _GEN_21020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21022 = 9'h2a == r_count_52_io_out ? io_r_42_b : _GEN_21021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21023 = 9'h2b == r_count_52_io_out ? io_r_43_b : _GEN_21022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21024 = 9'h2c == r_count_52_io_out ? io_r_44_b : _GEN_21023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21025 = 9'h2d == r_count_52_io_out ? io_r_45_b : _GEN_21024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21026 = 9'h2e == r_count_52_io_out ? io_r_46_b : _GEN_21025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21027 = 9'h2f == r_count_52_io_out ? io_r_47_b : _GEN_21026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21028 = 9'h30 == r_count_52_io_out ? io_r_48_b : _GEN_21027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21029 = 9'h31 == r_count_52_io_out ? io_r_49_b : _GEN_21028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21030 = 9'h32 == r_count_52_io_out ? io_r_50_b : _GEN_21029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21031 = 9'h33 == r_count_52_io_out ? io_r_51_b : _GEN_21030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21032 = 9'h34 == r_count_52_io_out ? io_r_52_b : _GEN_21031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21033 = 9'h35 == r_count_52_io_out ? io_r_53_b : _GEN_21032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21034 = 9'h36 == r_count_52_io_out ? io_r_54_b : _GEN_21033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21035 = 9'h37 == r_count_52_io_out ? io_r_55_b : _GEN_21034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21036 = 9'h38 == r_count_52_io_out ? io_r_56_b : _GEN_21035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21037 = 9'h39 == r_count_52_io_out ? io_r_57_b : _GEN_21036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21038 = 9'h3a == r_count_52_io_out ? io_r_58_b : _GEN_21037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21039 = 9'h3b == r_count_52_io_out ? io_r_59_b : _GEN_21038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21040 = 9'h3c == r_count_52_io_out ? io_r_60_b : _GEN_21039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21041 = 9'h3d == r_count_52_io_out ? io_r_61_b : _GEN_21040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21042 = 9'h3e == r_count_52_io_out ? io_r_62_b : _GEN_21041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21043 = 9'h3f == r_count_52_io_out ? io_r_63_b : _GEN_21042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21044 = 9'h40 == r_count_52_io_out ? io_r_64_b : _GEN_21043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21045 = 9'h41 == r_count_52_io_out ? io_r_65_b : _GEN_21044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21046 = 9'h42 == r_count_52_io_out ? io_r_66_b : _GEN_21045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21047 = 9'h43 == r_count_52_io_out ? io_r_67_b : _GEN_21046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21048 = 9'h44 == r_count_52_io_out ? io_r_68_b : _GEN_21047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21049 = 9'h45 == r_count_52_io_out ? io_r_69_b : _GEN_21048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21050 = 9'h46 == r_count_52_io_out ? io_r_70_b : _GEN_21049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21051 = 9'h47 == r_count_52_io_out ? io_r_71_b : _GEN_21050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21052 = 9'h48 == r_count_52_io_out ? io_r_72_b : _GEN_21051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21053 = 9'h49 == r_count_52_io_out ? io_r_73_b : _GEN_21052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21054 = 9'h4a == r_count_52_io_out ? io_r_74_b : _GEN_21053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21055 = 9'h4b == r_count_52_io_out ? io_r_75_b : _GEN_21054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21056 = 9'h4c == r_count_52_io_out ? io_r_76_b : _GEN_21055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21057 = 9'h4d == r_count_52_io_out ? io_r_77_b : _GEN_21056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21058 = 9'h4e == r_count_52_io_out ? io_r_78_b : _GEN_21057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21059 = 9'h4f == r_count_52_io_out ? io_r_79_b : _GEN_21058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21060 = 9'h50 == r_count_52_io_out ? io_r_80_b : _GEN_21059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21061 = 9'h51 == r_count_52_io_out ? io_r_81_b : _GEN_21060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21062 = 9'h52 == r_count_52_io_out ? io_r_82_b : _GEN_21061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21063 = 9'h53 == r_count_52_io_out ? io_r_83_b : _GEN_21062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21064 = 9'h54 == r_count_52_io_out ? io_r_84_b : _GEN_21063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21065 = 9'h55 == r_count_52_io_out ? io_r_85_b : _GEN_21064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21066 = 9'h56 == r_count_52_io_out ? io_r_86_b : _GEN_21065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21067 = 9'h57 == r_count_52_io_out ? io_r_87_b : _GEN_21066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21068 = 9'h58 == r_count_52_io_out ? io_r_88_b : _GEN_21067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21069 = 9'h59 == r_count_52_io_out ? io_r_89_b : _GEN_21068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21070 = 9'h5a == r_count_52_io_out ? io_r_90_b : _GEN_21069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21071 = 9'h5b == r_count_52_io_out ? io_r_91_b : _GEN_21070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21072 = 9'h5c == r_count_52_io_out ? io_r_92_b : _GEN_21071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21073 = 9'h5d == r_count_52_io_out ? io_r_93_b : _GEN_21072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21074 = 9'h5e == r_count_52_io_out ? io_r_94_b : _GEN_21073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21075 = 9'h5f == r_count_52_io_out ? io_r_95_b : _GEN_21074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21076 = 9'h60 == r_count_52_io_out ? io_r_96_b : _GEN_21075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21077 = 9'h61 == r_count_52_io_out ? io_r_97_b : _GEN_21076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21078 = 9'h62 == r_count_52_io_out ? io_r_98_b : _GEN_21077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21079 = 9'h63 == r_count_52_io_out ? io_r_99_b : _GEN_21078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21080 = 9'h64 == r_count_52_io_out ? io_r_100_b : _GEN_21079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21081 = 9'h65 == r_count_52_io_out ? io_r_101_b : _GEN_21080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21082 = 9'h66 == r_count_52_io_out ? io_r_102_b : _GEN_21081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21083 = 9'h67 == r_count_52_io_out ? io_r_103_b : _GEN_21082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21084 = 9'h68 == r_count_52_io_out ? io_r_104_b : _GEN_21083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21085 = 9'h69 == r_count_52_io_out ? io_r_105_b : _GEN_21084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21086 = 9'h6a == r_count_52_io_out ? io_r_106_b : _GEN_21085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21087 = 9'h6b == r_count_52_io_out ? io_r_107_b : _GEN_21086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21088 = 9'h6c == r_count_52_io_out ? io_r_108_b : _GEN_21087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21089 = 9'h6d == r_count_52_io_out ? io_r_109_b : _GEN_21088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21090 = 9'h6e == r_count_52_io_out ? io_r_110_b : _GEN_21089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21091 = 9'h6f == r_count_52_io_out ? io_r_111_b : _GEN_21090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21092 = 9'h70 == r_count_52_io_out ? io_r_112_b : _GEN_21091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21093 = 9'h71 == r_count_52_io_out ? io_r_113_b : _GEN_21092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21094 = 9'h72 == r_count_52_io_out ? io_r_114_b : _GEN_21093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21095 = 9'h73 == r_count_52_io_out ? io_r_115_b : _GEN_21094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21096 = 9'h74 == r_count_52_io_out ? io_r_116_b : _GEN_21095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21097 = 9'h75 == r_count_52_io_out ? io_r_117_b : _GEN_21096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21098 = 9'h76 == r_count_52_io_out ? io_r_118_b : _GEN_21097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21099 = 9'h77 == r_count_52_io_out ? io_r_119_b : _GEN_21098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21100 = 9'h78 == r_count_52_io_out ? io_r_120_b : _GEN_21099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21101 = 9'h79 == r_count_52_io_out ? io_r_121_b : _GEN_21100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21102 = 9'h7a == r_count_52_io_out ? io_r_122_b : _GEN_21101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21103 = 9'h7b == r_count_52_io_out ? io_r_123_b : _GEN_21102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21104 = 9'h7c == r_count_52_io_out ? io_r_124_b : _GEN_21103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21105 = 9'h7d == r_count_52_io_out ? io_r_125_b : _GEN_21104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21106 = 9'h7e == r_count_52_io_out ? io_r_126_b : _GEN_21105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21107 = 9'h7f == r_count_52_io_out ? io_r_127_b : _GEN_21106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21108 = 9'h80 == r_count_52_io_out ? io_r_128_b : _GEN_21107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21109 = 9'h81 == r_count_52_io_out ? io_r_129_b : _GEN_21108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21110 = 9'h82 == r_count_52_io_out ? io_r_130_b : _GEN_21109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21111 = 9'h83 == r_count_52_io_out ? io_r_131_b : _GEN_21110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21112 = 9'h84 == r_count_52_io_out ? io_r_132_b : _GEN_21111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21113 = 9'h85 == r_count_52_io_out ? io_r_133_b : _GEN_21112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21114 = 9'h86 == r_count_52_io_out ? io_r_134_b : _GEN_21113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21115 = 9'h87 == r_count_52_io_out ? io_r_135_b : _GEN_21114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21116 = 9'h88 == r_count_52_io_out ? io_r_136_b : _GEN_21115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21117 = 9'h89 == r_count_52_io_out ? io_r_137_b : _GEN_21116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21118 = 9'h8a == r_count_52_io_out ? io_r_138_b : _GEN_21117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21119 = 9'h8b == r_count_52_io_out ? io_r_139_b : _GEN_21118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21120 = 9'h8c == r_count_52_io_out ? io_r_140_b : _GEN_21119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21121 = 9'h8d == r_count_52_io_out ? io_r_141_b : _GEN_21120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21122 = 9'h8e == r_count_52_io_out ? io_r_142_b : _GEN_21121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21123 = 9'h8f == r_count_52_io_out ? io_r_143_b : _GEN_21122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21124 = 9'h90 == r_count_52_io_out ? io_r_144_b : _GEN_21123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21125 = 9'h91 == r_count_52_io_out ? io_r_145_b : _GEN_21124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21126 = 9'h92 == r_count_52_io_out ? io_r_146_b : _GEN_21125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21127 = 9'h93 == r_count_52_io_out ? io_r_147_b : _GEN_21126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21128 = 9'h94 == r_count_52_io_out ? io_r_148_b : _GEN_21127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21129 = 9'h95 == r_count_52_io_out ? io_r_149_b : _GEN_21128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21130 = 9'h96 == r_count_52_io_out ? io_r_150_b : _GEN_21129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21131 = 9'h97 == r_count_52_io_out ? io_r_151_b : _GEN_21130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21132 = 9'h98 == r_count_52_io_out ? io_r_152_b : _GEN_21131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21133 = 9'h99 == r_count_52_io_out ? io_r_153_b : _GEN_21132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21134 = 9'h9a == r_count_52_io_out ? io_r_154_b : _GEN_21133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21135 = 9'h9b == r_count_52_io_out ? io_r_155_b : _GEN_21134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21136 = 9'h9c == r_count_52_io_out ? io_r_156_b : _GEN_21135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21137 = 9'h9d == r_count_52_io_out ? io_r_157_b : _GEN_21136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21138 = 9'h9e == r_count_52_io_out ? io_r_158_b : _GEN_21137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21139 = 9'h9f == r_count_52_io_out ? io_r_159_b : _GEN_21138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21140 = 9'ha0 == r_count_52_io_out ? io_r_160_b : _GEN_21139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21141 = 9'ha1 == r_count_52_io_out ? io_r_161_b : _GEN_21140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21142 = 9'ha2 == r_count_52_io_out ? io_r_162_b : _GEN_21141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21143 = 9'ha3 == r_count_52_io_out ? io_r_163_b : _GEN_21142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21144 = 9'ha4 == r_count_52_io_out ? io_r_164_b : _GEN_21143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21145 = 9'ha5 == r_count_52_io_out ? io_r_165_b : _GEN_21144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21146 = 9'ha6 == r_count_52_io_out ? io_r_166_b : _GEN_21145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21147 = 9'ha7 == r_count_52_io_out ? io_r_167_b : _GEN_21146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21148 = 9'ha8 == r_count_52_io_out ? io_r_168_b : _GEN_21147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21149 = 9'ha9 == r_count_52_io_out ? io_r_169_b : _GEN_21148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21150 = 9'haa == r_count_52_io_out ? io_r_170_b : _GEN_21149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21151 = 9'hab == r_count_52_io_out ? io_r_171_b : _GEN_21150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21152 = 9'hac == r_count_52_io_out ? io_r_172_b : _GEN_21151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21153 = 9'had == r_count_52_io_out ? io_r_173_b : _GEN_21152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21154 = 9'hae == r_count_52_io_out ? io_r_174_b : _GEN_21153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21155 = 9'haf == r_count_52_io_out ? io_r_175_b : _GEN_21154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21156 = 9'hb0 == r_count_52_io_out ? io_r_176_b : _GEN_21155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21157 = 9'hb1 == r_count_52_io_out ? io_r_177_b : _GEN_21156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21158 = 9'hb2 == r_count_52_io_out ? io_r_178_b : _GEN_21157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21159 = 9'hb3 == r_count_52_io_out ? io_r_179_b : _GEN_21158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21160 = 9'hb4 == r_count_52_io_out ? io_r_180_b : _GEN_21159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21161 = 9'hb5 == r_count_52_io_out ? io_r_181_b : _GEN_21160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21162 = 9'hb6 == r_count_52_io_out ? io_r_182_b : _GEN_21161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21163 = 9'hb7 == r_count_52_io_out ? io_r_183_b : _GEN_21162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21164 = 9'hb8 == r_count_52_io_out ? io_r_184_b : _GEN_21163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21165 = 9'hb9 == r_count_52_io_out ? io_r_185_b : _GEN_21164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21166 = 9'hba == r_count_52_io_out ? io_r_186_b : _GEN_21165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21167 = 9'hbb == r_count_52_io_out ? io_r_187_b : _GEN_21166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21168 = 9'hbc == r_count_52_io_out ? io_r_188_b : _GEN_21167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21169 = 9'hbd == r_count_52_io_out ? io_r_189_b : _GEN_21168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21170 = 9'hbe == r_count_52_io_out ? io_r_190_b : _GEN_21169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21171 = 9'hbf == r_count_52_io_out ? io_r_191_b : _GEN_21170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21172 = 9'hc0 == r_count_52_io_out ? io_r_192_b : _GEN_21171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21173 = 9'hc1 == r_count_52_io_out ? io_r_193_b : _GEN_21172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21174 = 9'hc2 == r_count_52_io_out ? io_r_194_b : _GEN_21173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21175 = 9'hc3 == r_count_52_io_out ? io_r_195_b : _GEN_21174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21176 = 9'hc4 == r_count_52_io_out ? io_r_196_b : _GEN_21175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21177 = 9'hc5 == r_count_52_io_out ? io_r_197_b : _GEN_21176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21178 = 9'hc6 == r_count_52_io_out ? io_r_198_b : _GEN_21177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21179 = 9'hc7 == r_count_52_io_out ? io_r_199_b : _GEN_21178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21180 = 9'hc8 == r_count_52_io_out ? io_r_200_b : _GEN_21179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21181 = 9'hc9 == r_count_52_io_out ? io_r_201_b : _GEN_21180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21182 = 9'hca == r_count_52_io_out ? io_r_202_b : _GEN_21181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21183 = 9'hcb == r_count_52_io_out ? io_r_203_b : _GEN_21182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21184 = 9'hcc == r_count_52_io_out ? io_r_204_b : _GEN_21183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21185 = 9'hcd == r_count_52_io_out ? io_r_205_b : _GEN_21184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21186 = 9'hce == r_count_52_io_out ? io_r_206_b : _GEN_21185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21187 = 9'hcf == r_count_52_io_out ? io_r_207_b : _GEN_21186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21188 = 9'hd0 == r_count_52_io_out ? io_r_208_b : _GEN_21187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21189 = 9'hd1 == r_count_52_io_out ? io_r_209_b : _GEN_21188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21190 = 9'hd2 == r_count_52_io_out ? io_r_210_b : _GEN_21189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21191 = 9'hd3 == r_count_52_io_out ? io_r_211_b : _GEN_21190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21192 = 9'hd4 == r_count_52_io_out ? io_r_212_b : _GEN_21191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21193 = 9'hd5 == r_count_52_io_out ? io_r_213_b : _GEN_21192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21194 = 9'hd6 == r_count_52_io_out ? io_r_214_b : _GEN_21193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21195 = 9'hd7 == r_count_52_io_out ? io_r_215_b : _GEN_21194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21196 = 9'hd8 == r_count_52_io_out ? io_r_216_b : _GEN_21195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21197 = 9'hd9 == r_count_52_io_out ? io_r_217_b : _GEN_21196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21198 = 9'hda == r_count_52_io_out ? io_r_218_b : _GEN_21197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21199 = 9'hdb == r_count_52_io_out ? io_r_219_b : _GEN_21198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21200 = 9'hdc == r_count_52_io_out ? io_r_220_b : _GEN_21199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21201 = 9'hdd == r_count_52_io_out ? io_r_221_b : _GEN_21200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21202 = 9'hde == r_count_52_io_out ? io_r_222_b : _GEN_21201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21203 = 9'hdf == r_count_52_io_out ? io_r_223_b : _GEN_21202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21204 = 9'he0 == r_count_52_io_out ? io_r_224_b : _GEN_21203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21205 = 9'he1 == r_count_52_io_out ? io_r_225_b : _GEN_21204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21206 = 9'he2 == r_count_52_io_out ? io_r_226_b : _GEN_21205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21207 = 9'he3 == r_count_52_io_out ? io_r_227_b : _GEN_21206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21208 = 9'he4 == r_count_52_io_out ? io_r_228_b : _GEN_21207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21209 = 9'he5 == r_count_52_io_out ? io_r_229_b : _GEN_21208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21210 = 9'he6 == r_count_52_io_out ? io_r_230_b : _GEN_21209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21211 = 9'he7 == r_count_52_io_out ? io_r_231_b : _GEN_21210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21212 = 9'he8 == r_count_52_io_out ? io_r_232_b : _GEN_21211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21213 = 9'he9 == r_count_52_io_out ? io_r_233_b : _GEN_21212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21214 = 9'hea == r_count_52_io_out ? io_r_234_b : _GEN_21213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21215 = 9'heb == r_count_52_io_out ? io_r_235_b : _GEN_21214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21216 = 9'hec == r_count_52_io_out ? io_r_236_b : _GEN_21215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21217 = 9'hed == r_count_52_io_out ? io_r_237_b : _GEN_21216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21218 = 9'hee == r_count_52_io_out ? io_r_238_b : _GEN_21217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21219 = 9'hef == r_count_52_io_out ? io_r_239_b : _GEN_21218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21220 = 9'hf0 == r_count_52_io_out ? io_r_240_b : _GEN_21219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21221 = 9'hf1 == r_count_52_io_out ? io_r_241_b : _GEN_21220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21222 = 9'hf2 == r_count_52_io_out ? io_r_242_b : _GEN_21221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21223 = 9'hf3 == r_count_52_io_out ? io_r_243_b : _GEN_21222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21224 = 9'hf4 == r_count_52_io_out ? io_r_244_b : _GEN_21223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21225 = 9'hf5 == r_count_52_io_out ? io_r_245_b : _GEN_21224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21226 = 9'hf6 == r_count_52_io_out ? io_r_246_b : _GEN_21225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21227 = 9'hf7 == r_count_52_io_out ? io_r_247_b : _GEN_21226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21228 = 9'hf8 == r_count_52_io_out ? io_r_248_b : _GEN_21227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21229 = 9'hf9 == r_count_52_io_out ? io_r_249_b : _GEN_21228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21230 = 9'hfa == r_count_52_io_out ? io_r_250_b : _GEN_21229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21231 = 9'hfb == r_count_52_io_out ? io_r_251_b : _GEN_21230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21232 = 9'hfc == r_count_52_io_out ? io_r_252_b : _GEN_21231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21233 = 9'hfd == r_count_52_io_out ? io_r_253_b : _GEN_21232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21234 = 9'hfe == r_count_52_io_out ? io_r_254_b : _GEN_21233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21235 = 9'hff == r_count_52_io_out ? io_r_255_b : _GEN_21234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21236 = 9'h100 == r_count_52_io_out ? io_r_256_b : _GEN_21235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21237 = 9'h101 == r_count_52_io_out ? io_r_257_b : _GEN_21236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21238 = 9'h102 == r_count_52_io_out ? io_r_258_b : _GEN_21237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21239 = 9'h103 == r_count_52_io_out ? io_r_259_b : _GEN_21238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21240 = 9'h104 == r_count_52_io_out ? io_r_260_b : _GEN_21239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21241 = 9'h105 == r_count_52_io_out ? io_r_261_b : _GEN_21240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21242 = 9'h106 == r_count_52_io_out ? io_r_262_b : _GEN_21241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21243 = 9'h107 == r_count_52_io_out ? io_r_263_b : _GEN_21242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21244 = 9'h108 == r_count_52_io_out ? io_r_264_b : _GEN_21243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21245 = 9'h109 == r_count_52_io_out ? io_r_265_b : _GEN_21244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21246 = 9'h10a == r_count_52_io_out ? io_r_266_b : _GEN_21245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21247 = 9'h10b == r_count_52_io_out ? io_r_267_b : _GEN_21246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21248 = 9'h10c == r_count_52_io_out ? io_r_268_b : _GEN_21247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21249 = 9'h10d == r_count_52_io_out ? io_r_269_b : _GEN_21248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21250 = 9'h10e == r_count_52_io_out ? io_r_270_b : _GEN_21249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21251 = 9'h10f == r_count_52_io_out ? io_r_271_b : _GEN_21250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21252 = 9'h110 == r_count_52_io_out ? io_r_272_b : _GEN_21251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21253 = 9'h111 == r_count_52_io_out ? io_r_273_b : _GEN_21252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21254 = 9'h112 == r_count_52_io_out ? io_r_274_b : _GEN_21253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21255 = 9'h113 == r_count_52_io_out ? io_r_275_b : _GEN_21254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21256 = 9'h114 == r_count_52_io_out ? io_r_276_b : _GEN_21255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21257 = 9'h115 == r_count_52_io_out ? io_r_277_b : _GEN_21256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21258 = 9'h116 == r_count_52_io_out ? io_r_278_b : _GEN_21257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21259 = 9'h117 == r_count_52_io_out ? io_r_279_b : _GEN_21258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21260 = 9'h118 == r_count_52_io_out ? io_r_280_b : _GEN_21259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21261 = 9'h119 == r_count_52_io_out ? io_r_281_b : _GEN_21260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21262 = 9'h11a == r_count_52_io_out ? io_r_282_b : _GEN_21261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21263 = 9'h11b == r_count_52_io_out ? io_r_283_b : _GEN_21262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21264 = 9'h11c == r_count_52_io_out ? io_r_284_b : _GEN_21263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21265 = 9'h11d == r_count_52_io_out ? io_r_285_b : _GEN_21264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21266 = 9'h11e == r_count_52_io_out ? io_r_286_b : _GEN_21265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21267 = 9'h11f == r_count_52_io_out ? io_r_287_b : _GEN_21266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21268 = 9'h120 == r_count_52_io_out ? io_r_288_b : _GEN_21267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21269 = 9'h121 == r_count_52_io_out ? io_r_289_b : _GEN_21268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21270 = 9'h122 == r_count_52_io_out ? io_r_290_b : _GEN_21269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21271 = 9'h123 == r_count_52_io_out ? io_r_291_b : _GEN_21270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21272 = 9'h124 == r_count_52_io_out ? io_r_292_b : _GEN_21271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21273 = 9'h125 == r_count_52_io_out ? io_r_293_b : _GEN_21272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21274 = 9'h126 == r_count_52_io_out ? io_r_294_b : _GEN_21273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21275 = 9'h127 == r_count_52_io_out ? io_r_295_b : _GEN_21274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21276 = 9'h128 == r_count_52_io_out ? io_r_296_b : _GEN_21275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21277 = 9'h129 == r_count_52_io_out ? io_r_297_b : _GEN_21276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21278 = 9'h12a == r_count_52_io_out ? io_r_298_b : _GEN_21277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21279 = 9'h12b == r_count_52_io_out ? io_r_299_b : _GEN_21278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21280 = 9'h12c == r_count_52_io_out ? io_r_300_b : _GEN_21279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21281 = 9'h12d == r_count_52_io_out ? io_r_301_b : _GEN_21280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21282 = 9'h12e == r_count_52_io_out ? io_r_302_b : _GEN_21281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21283 = 9'h12f == r_count_52_io_out ? io_r_303_b : _GEN_21282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21284 = 9'h130 == r_count_52_io_out ? io_r_304_b : _GEN_21283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21285 = 9'h131 == r_count_52_io_out ? io_r_305_b : _GEN_21284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21286 = 9'h132 == r_count_52_io_out ? io_r_306_b : _GEN_21285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21287 = 9'h133 == r_count_52_io_out ? io_r_307_b : _GEN_21286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21288 = 9'h134 == r_count_52_io_out ? io_r_308_b : _GEN_21287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21289 = 9'h135 == r_count_52_io_out ? io_r_309_b : _GEN_21288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21290 = 9'h136 == r_count_52_io_out ? io_r_310_b : _GEN_21289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21291 = 9'h137 == r_count_52_io_out ? io_r_311_b : _GEN_21290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21292 = 9'h138 == r_count_52_io_out ? io_r_312_b : _GEN_21291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21293 = 9'h139 == r_count_52_io_out ? io_r_313_b : _GEN_21292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21294 = 9'h13a == r_count_52_io_out ? io_r_314_b : _GEN_21293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21295 = 9'h13b == r_count_52_io_out ? io_r_315_b : _GEN_21294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21296 = 9'h13c == r_count_52_io_out ? io_r_316_b : _GEN_21295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21297 = 9'h13d == r_count_52_io_out ? io_r_317_b : _GEN_21296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21298 = 9'h13e == r_count_52_io_out ? io_r_318_b : _GEN_21297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21299 = 9'h13f == r_count_52_io_out ? io_r_319_b : _GEN_21298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21300 = 9'h140 == r_count_52_io_out ? io_r_320_b : _GEN_21299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21301 = 9'h141 == r_count_52_io_out ? io_r_321_b : _GEN_21300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21302 = 9'h142 == r_count_52_io_out ? io_r_322_b : _GEN_21301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21303 = 9'h143 == r_count_52_io_out ? io_r_323_b : _GEN_21302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21304 = 9'h144 == r_count_52_io_out ? io_r_324_b : _GEN_21303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21305 = 9'h145 == r_count_52_io_out ? io_r_325_b : _GEN_21304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21306 = 9'h146 == r_count_52_io_out ? io_r_326_b : _GEN_21305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21307 = 9'h147 == r_count_52_io_out ? io_r_327_b : _GEN_21306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21308 = 9'h148 == r_count_52_io_out ? io_r_328_b : _GEN_21307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21309 = 9'h149 == r_count_52_io_out ? io_r_329_b : _GEN_21308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21310 = 9'h14a == r_count_52_io_out ? io_r_330_b : _GEN_21309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21311 = 9'h14b == r_count_52_io_out ? io_r_331_b : _GEN_21310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21312 = 9'h14c == r_count_52_io_out ? io_r_332_b : _GEN_21311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21313 = 9'h14d == r_count_52_io_out ? io_r_333_b : _GEN_21312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21314 = 9'h14e == r_count_52_io_out ? io_r_334_b : _GEN_21313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21315 = 9'h14f == r_count_52_io_out ? io_r_335_b : _GEN_21314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21316 = 9'h150 == r_count_52_io_out ? io_r_336_b : _GEN_21315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21317 = 9'h151 == r_count_52_io_out ? io_r_337_b : _GEN_21316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21318 = 9'h152 == r_count_52_io_out ? io_r_338_b : _GEN_21317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21319 = 9'h153 == r_count_52_io_out ? io_r_339_b : _GEN_21318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21320 = 9'h154 == r_count_52_io_out ? io_r_340_b : _GEN_21319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21321 = 9'h155 == r_count_52_io_out ? io_r_341_b : _GEN_21320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21322 = 9'h156 == r_count_52_io_out ? io_r_342_b : _GEN_21321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21323 = 9'h157 == r_count_52_io_out ? io_r_343_b : _GEN_21322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21324 = 9'h158 == r_count_52_io_out ? io_r_344_b : _GEN_21323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21325 = 9'h159 == r_count_52_io_out ? io_r_345_b : _GEN_21324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21326 = 9'h15a == r_count_52_io_out ? io_r_346_b : _GEN_21325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21327 = 9'h15b == r_count_52_io_out ? io_r_347_b : _GEN_21326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21328 = 9'h15c == r_count_52_io_out ? io_r_348_b : _GEN_21327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21329 = 9'h15d == r_count_52_io_out ? io_r_349_b : _GEN_21328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21330 = 9'h15e == r_count_52_io_out ? io_r_350_b : _GEN_21329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21331 = 9'h15f == r_count_52_io_out ? io_r_351_b : _GEN_21330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21332 = 9'h160 == r_count_52_io_out ? io_r_352_b : _GEN_21331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21333 = 9'h161 == r_count_52_io_out ? io_r_353_b : _GEN_21332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21334 = 9'h162 == r_count_52_io_out ? io_r_354_b : _GEN_21333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21335 = 9'h163 == r_count_52_io_out ? io_r_355_b : _GEN_21334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21336 = 9'h164 == r_count_52_io_out ? io_r_356_b : _GEN_21335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21337 = 9'h165 == r_count_52_io_out ? io_r_357_b : _GEN_21336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21338 = 9'h166 == r_count_52_io_out ? io_r_358_b : _GEN_21337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21339 = 9'h167 == r_count_52_io_out ? io_r_359_b : _GEN_21338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21340 = 9'h168 == r_count_52_io_out ? io_r_360_b : _GEN_21339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21341 = 9'h169 == r_count_52_io_out ? io_r_361_b : _GEN_21340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21342 = 9'h16a == r_count_52_io_out ? io_r_362_b : _GEN_21341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21343 = 9'h16b == r_count_52_io_out ? io_r_363_b : _GEN_21342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21344 = 9'h16c == r_count_52_io_out ? io_r_364_b : _GEN_21343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21345 = 9'h16d == r_count_52_io_out ? io_r_365_b : _GEN_21344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21346 = 9'h16e == r_count_52_io_out ? io_r_366_b : _GEN_21345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21347 = 9'h16f == r_count_52_io_out ? io_r_367_b : _GEN_21346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21348 = 9'h170 == r_count_52_io_out ? io_r_368_b : _GEN_21347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21349 = 9'h171 == r_count_52_io_out ? io_r_369_b : _GEN_21348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21350 = 9'h172 == r_count_52_io_out ? io_r_370_b : _GEN_21349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21351 = 9'h173 == r_count_52_io_out ? io_r_371_b : _GEN_21350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21352 = 9'h174 == r_count_52_io_out ? io_r_372_b : _GEN_21351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21353 = 9'h175 == r_count_52_io_out ? io_r_373_b : _GEN_21352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21354 = 9'h176 == r_count_52_io_out ? io_r_374_b : _GEN_21353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21355 = 9'h177 == r_count_52_io_out ? io_r_375_b : _GEN_21354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21356 = 9'h178 == r_count_52_io_out ? io_r_376_b : _GEN_21355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21357 = 9'h179 == r_count_52_io_out ? io_r_377_b : _GEN_21356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21358 = 9'h17a == r_count_52_io_out ? io_r_378_b : _GEN_21357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21359 = 9'h17b == r_count_52_io_out ? io_r_379_b : _GEN_21358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21360 = 9'h17c == r_count_52_io_out ? io_r_380_b : _GEN_21359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21361 = 9'h17d == r_count_52_io_out ? io_r_381_b : _GEN_21360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21362 = 9'h17e == r_count_52_io_out ? io_r_382_b : _GEN_21361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21363 = 9'h17f == r_count_52_io_out ? io_r_383_b : _GEN_21362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21364 = 9'h180 == r_count_52_io_out ? io_r_384_b : _GEN_21363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21365 = 9'h181 == r_count_52_io_out ? io_r_385_b : _GEN_21364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21366 = 9'h182 == r_count_52_io_out ? io_r_386_b : _GEN_21365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21367 = 9'h183 == r_count_52_io_out ? io_r_387_b : _GEN_21366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21368 = 9'h184 == r_count_52_io_out ? io_r_388_b : _GEN_21367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21369 = 9'h185 == r_count_52_io_out ? io_r_389_b : _GEN_21368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21370 = 9'h186 == r_count_52_io_out ? io_r_390_b : _GEN_21369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21371 = 9'h187 == r_count_52_io_out ? io_r_391_b : _GEN_21370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21372 = 9'h188 == r_count_52_io_out ? io_r_392_b : _GEN_21371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21373 = 9'h189 == r_count_52_io_out ? io_r_393_b : _GEN_21372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21374 = 9'h18a == r_count_52_io_out ? io_r_394_b : _GEN_21373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21375 = 9'h18b == r_count_52_io_out ? io_r_395_b : _GEN_21374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21376 = 9'h18c == r_count_52_io_out ? io_r_396_b : _GEN_21375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21377 = 9'h18d == r_count_52_io_out ? io_r_397_b : _GEN_21376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21378 = 9'h18e == r_count_52_io_out ? io_r_398_b : _GEN_21377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21381 = 9'h1 == r_count_53_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21382 = 9'h2 == r_count_53_io_out ? io_r_2_b : _GEN_21381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21383 = 9'h3 == r_count_53_io_out ? io_r_3_b : _GEN_21382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21384 = 9'h4 == r_count_53_io_out ? io_r_4_b : _GEN_21383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21385 = 9'h5 == r_count_53_io_out ? io_r_5_b : _GEN_21384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21386 = 9'h6 == r_count_53_io_out ? io_r_6_b : _GEN_21385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21387 = 9'h7 == r_count_53_io_out ? io_r_7_b : _GEN_21386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21388 = 9'h8 == r_count_53_io_out ? io_r_8_b : _GEN_21387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21389 = 9'h9 == r_count_53_io_out ? io_r_9_b : _GEN_21388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21390 = 9'ha == r_count_53_io_out ? io_r_10_b : _GEN_21389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21391 = 9'hb == r_count_53_io_out ? io_r_11_b : _GEN_21390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21392 = 9'hc == r_count_53_io_out ? io_r_12_b : _GEN_21391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21393 = 9'hd == r_count_53_io_out ? io_r_13_b : _GEN_21392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21394 = 9'he == r_count_53_io_out ? io_r_14_b : _GEN_21393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21395 = 9'hf == r_count_53_io_out ? io_r_15_b : _GEN_21394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21396 = 9'h10 == r_count_53_io_out ? io_r_16_b : _GEN_21395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21397 = 9'h11 == r_count_53_io_out ? io_r_17_b : _GEN_21396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21398 = 9'h12 == r_count_53_io_out ? io_r_18_b : _GEN_21397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21399 = 9'h13 == r_count_53_io_out ? io_r_19_b : _GEN_21398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21400 = 9'h14 == r_count_53_io_out ? io_r_20_b : _GEN_21399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21401 = 9'h15 == r_count_53_io_out ? io_r_21_b : _GEN_21400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21402 = 9'h16 == r_count_53_io_out ? io_r_22_b : _GEN_21401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21403 = 9'h17 == r_count_53_io_out ? io_r_23_b : _GEN_21402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21404 = 9'h18 == r_count_53_io_out ? io_r_24_b : _GEN_21403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21405 = 9'h19 == r_count_53_io_out ? io_r_25_b : _GEN_21404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21406 = 9'h1a == r_count_53_io_out ? io_r_26_b : _GEN_21405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21407 = 9'h1b == r_count_53_io_out ? io_r_27_b : _GEN_21406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21408 = 9'h1c == r_count_53_io_out ? io_r_28_b : _GEN_21407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21409 = 9'h1d == r_count_53_io_out ? io_r_29_b : _GEN_21408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21410 = 9'h1e == r_count_53_io_out ? io_r_30_b : _GEN_21409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21411 = 9'h1f == r_count_53_io_out ? io_r_31_b : _GEN_21410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21412 = 9'h20 == r_count_53_io_out ? io_r_32_b : _GEN_21411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21413 = 9'h21 == r_count_53_io_out ? io_r_33_b : _GEN_21412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21414 = 9'h22 == r_count_53_io_out ? io_r_34_b : _GEN_21413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21415 = 9'h23 == r_count_53_io_out ? io_r_35_b : _GEN_21414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21416 = 9'h24 == r_count_53_io_out ? io_r_36_b : _GEN_21415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21417 = 9'h25 == r_count_53_io_out ? io_r_37_b : _GEN_21416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21418 = 9'h26 == r_count_53_io_out ? io_r_38_b : _GEN_21417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21419 = 9'h27 == r_count_53_io_out ? io_r_39_b : _GEN_21418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21420 = 9'h28 == r_count_53_io_out ? io_r_40_b : _GEN_21419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21421 = 9'h29 == r_count_53_io_out ? io_r_41_b : _GEN_21420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21422 = 9'h2a == r_count_53_io_out ? io_r_42_b : _GEN_21421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21423 = 9'h2b == r_count_53_io_out ? io_r_43_b : _GEN_21422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21424 = 9'h2c == r_count_53_io_out ? io_r_44_b : _GEN_21423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21425 = 9'h2d == r_count_53_io_out ? io_r_45_b : _GEN_21424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21426 = 9'h2e == r_count_53_io_out ? io_r_46_b : _GEN_21425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21427 = 9'h2f == r_count_53_io_out ? io_r_47_b : _GEN_21426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21428 = 9'h30 == r_count_53_io_out ? io_r_48_b : _GEN_21427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21429 = 9'h31 == r_count_53_io_out ? io_r_49_b : _GEN_21428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21430 = 9'h32 == r_count_53_io_out ? io_r_50_b : _GEN_21429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21431 = 9'h33 == r_count_53_io_out ? io_r_51_b : _GEN_21430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21432 = 9'h34 == r_count_53_io_out ? io_r_52_b : _GEN_21431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21433 = 9'h35 == r_count_53_io_out ? io_r_53_b : _GEN_21432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21434 = 9'h36 == r_count_53_io_out ? io_r_54_b : _GEN_21433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21435 = 9'h37 == r_count_53_io_out ? io_r_55_b : _GEN_21434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21436 = 9'h38 == r_count_53_io_out ? io_r_56_b : _GEN_21435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21437 = 9'h39 == r_count_53_io_out ? io_r_57_b : _GEN_21436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21438 = 9'h3a == r_count_53_io_out ? io_r_58_b : _GEN_21437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21439 = 9'h3b == r_count_53_io_out ? io_r_59_b : _GEN_21438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21440 = 9'h3c == r_count_53_io_out ? io_r_60_b : _GEN_21439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21441 = 9'h3d == r_count_53_io_out ? io_r_61_b : _GEN_21440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21442 = 9'h3e == r_count_53_io_out ? io_r_62_b : _GEN_21441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21443 = 9'h3f == r_count_53_io_out ? io_r_63_b : _GEN_21442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21444 = 9'h40 == r_count_53_io_out ? io_r_64_b : _GEN_21443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21445 = 9'h41 == r_count_53_io_out ? io_r_65_b : _GEN_21444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21446 = 9'h42 == r_count_53_io_out ? io_r_66_b : _GEN_21445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21447 = 9'h43 == r_count_53_io_out ? io_r_67_b : _GEN_21446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21448 = 9'h44 == r_count_53_io_out ? io_r_68_b : _GEN_21447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21449 = 9'h45 == r_count_53_io_out ? io_r_69_b : _GEN_21448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21450 = 9'h46 == r_count_53_io_out ? io_r_70_b : _GEN_21449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21451 = 9'h47 == r_count_53_io_out ? io_r_71_b : _GEN_21450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21452 = 9'h48 == r_count_53_io_out ? io_r_72_b : _GEN_21451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21453 = 9'h49 == r_count_53_io_out ? io_r_73_b : _GEN_21452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21454 = 9'h4a == r_count_53_io_out ? io_r_74_b : _GEN_21453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21455 = 9'h4b == r_count_53_io_out ? io_r_75_b : _GEN_21454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21456 = 9'h4c == r_count_53_io_out ? io_r_76_b : _GEN_21455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21457 = 9'h4d == r_count_53_io_out ? io_r_77_b : _GEN_21456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21458 = 9'h4e == r_count_53_io_out ? io_r_78_b : _GEN_21457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21459 = 9'h4f == r_count_53_io_out ? io_r_79_b : _GEN_21458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21460 = 9'h50 == r_count_53_io_out ? io_r_80_b : _GEN_21459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21461 = 9'h51 == r_count_53_io_out ? io_r_81_b : _GEN_21460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21462 = 9'h52 == r_count_53_io_out ? io_r_82_b : _GEN_21461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21463 = 9'h53 == r_count_53_io_out ? io_r_83_b : _GEN_21462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21464 = 9'h54 == r_count_53_io_out ? io_r_84_b : _GEN_21463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21465 = 9'h55 == r_count_53_io_out ? io_r_85_b : _GEN_21464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21466 = 9'h56 == r_count_53_io_out ? io_r_86_b : _GEN_21465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21467 = 9'h57 == r_count_53_io_out ? io_r_87_b : _GEN_21466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21468 = 9'h58 == r_count_53_io_out ? io_r_88_b : _GEN_21467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21469 = 9'h59 == r_count_53_io_out ? io_r_89_b : _GEN_21468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21470 = 9'h5a == r_count_53_io_out ? io_r_90_b : _GEN_21469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21471 = 9'h5b == r_count_53_io_out ? io_r_91_b : _GEN_21470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21472 = 9'h5c == r_count_53_io_out ? io_r_92_b : _GEN_21471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21473 = 9'h5d == r_count_53_io_out ? io_r_93_b : _GEN_21472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21474 = 9'h5e == r_count_53_io_out ? io_r_94_b : _GEN_21473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21475 = 9'h5f == r_count_53_io_out ? io_r_95_b : _GEN_21474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21476 = 9'h60 == r_count_53_io_out ? io_r_96_b : _GEN_21475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21477 = 9'h61 == r_count_53_io_out ? io_r_97_b : _GEN_21476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21478 = 9'h62 == r_count_53_io_out ? io_r_98_b : _GEN_21477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21479 = 9'h63 == r_count_53_io_out ? io_r_99_b : _GEN_21478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21480 = 9'h64 == r_count_53_io_out ? io_r_100_b : _GEN_21479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21481 = 9'h65 == r_count_53_io_out ? io_r_101_b : _GEN_21480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21482 = 9'h66 == r_count_53_io_out ? io_r_102_b : _GEN_21481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21483 = 9'h67 == r_count_53_io_out ? io_r_103_b : _GEN_21482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21484 = 9'h68 == r_count_53_io_out ? io_r_104_b : _GEN_21483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21485 = 9'h69 == r_count_53_io_out ? io_r_105_b : _GEN_21484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21486 = 9'h6a == r_count_53_io_out ? io_r_106_b : _GEN_21485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21487 = 9'h6b == r_count_53_io_out ? io_r_107_b : _GEN_21486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21488 = 9'h6c == r_count_53_io_out ? io_r_108_b : _GEN_21487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21489 = 9'h6d == r_count_53_io_out ? io_r_109_b : _GEN_21488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21490 = 9'h6e == r_count_53_io_out ? io_r_110_b : _GEN_21489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21491 = 9'h6f == r_count_53_io_out ? io_r_111_b : _GEN_21490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21492 = 9'h70 == r_count_53_io_out ? io_r_112_b : _GEN_21491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21493 = 9'h71 == r_count_53_io_out ? io_r_113_b : _GEN_21492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21494 = 9'h72 == r_count_53_io_out ? io_r_114_b : _GEN_21493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21495 = 9'h73 == r_count_53_io_out ? io_r_115_b : _GEN_21494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21496 = 9'h74 == r_count_53_io_out ? io_r_116_b : _GEN_21495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21497 = 9'h75 == r_count_53_io_out ? io_r_117_b : _GEN_21496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21498 = 9'h76 == r_count_53_io_out ? io_r_118_b : _GEN_21497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21499 = 9'h77 == r_count_53_io_out ? io_r_119_b : _GEN_21498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21500 = 9'h78 == r_count_53_io_out ? io_r_120_b : _GEN_21499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21501 = 9'h79 == r_count_53_io_out ? io_r_121_b : _GEN_21500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21502 = 9'h7a == r_count_53_io_out ? io_r_122_b : _GEN_21501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21503 = 9'h7b == r_count_53_io_out ? io_r_123_b : _GEN_21502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21504 = 9'h7c == r_count_53_io_out ? io_r_124_b : _GEN_21503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21505 = 9'h7d == r_count_53_io_out ? io_r_125_b : _GEN_21504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21506 = 9'h7e == r_count_53_io_out ? io_r_126_b : _GEN_21505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21507 = 9'h7f == r_count_53_io_out ? io_r_127_b : _GEN_21506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21508 = 9'h80 == r_count_53_io_out ? io_r_128_b : _GEN_21507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21509 = 9'h81 == r_count_53_io_out ? io_r_129_b : _GEN_21508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21510 = 9'h82 == r_count_53_io_out ? io_r_130_b : _GEN_21509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21511 = 9'h83 == r_count_53_io_out ? io_r_131_b : _GEN_21510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21512 = 9'h84 == r_count_53_io_out ? io_r_132_b : _GEN_21511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21513 = 9'h85 == r_count_53_io_out ? io_r_133_b : _GEN_21512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21514 = 9'h86 == r_count_53_io_out ? io_r_134_b : _GEN_21513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21515 = 9'h87 == r_count_53_io_out ? io_r_135_b : _GEN_21514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21516 = 9'h88 == r_count_53_io_out ? io_r_136_b : _GEN_21515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21517 = 9'h89 == r_count_53_io_out ? io_r_137_b : _GEN_21516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21518 = 9'h8a == r_count_53_io_out ? io_r_138_b : _GEN_21517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21519 = 9'h8b == r_count_53_io_out ? io_r_139_b : _GEN_21518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21520 = 9'h8c == r_count_53_io_out ? io_r_140_b : _GEN_21519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21521 = 9'h8d == r_count_53_io_out ? io_r_141_b : _GEN_21520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21522 = 9'h8e == r_count_53_io_out ? io_r_142_b : _GEN_21521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21523 = 9'h8f == r_count_53_io_out ? io_r_143_b : _GEN_21522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21524 = 9'h90 == r_count_53_io_out ? io_r_144_b : _GEN_21523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21525 = 9'h91 == r_count_53_io_out ? io_r_145_b : _GEN_21524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21526 = 9'h92 == r_count_53_io_out ? io_r_146_b : _GEN_21525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21527 = 9'h93 == r_count_53_io_out ? io_r_147_b : _GEN_21526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21528 = 9'h94 == r_count_53_io_out ? io_r_148_b : _GEN_21527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21529 = 9'h95 == r_count_53_io_out ? io_r_149_b : _GEN_21528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21530 = 9'h96 == r_count_53_io_out ? io_r_150_b : _GEN_21529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21531 = 9'h97 == r_count_53_io_out ? io_r_151_b : _GEN_21530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21532 = 9'h98 == r_count_53_io_out ? io_r_152_b : _GEN_21531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21533 = 9'h99 == r_count_53_io_out ? io_r_153_b : _GEN_21532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21534 = 9'h9a == r_count_53_io_out ? io_r_154_b : _GEN_21533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21535 = 9'h9b == r_count_53_io_out ? io_r_155_b : _GEN_21534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21536 = 9'h9c == r_count_53_io_out ? io_r_156_b : _GEN_21535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21537 = 9'h9d == r_count_53_io_out ? io_r_157_b : _GEN_21536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21538 = 9'h9e == r_count_53_io_out ? io_r_158_b : _GEN_21537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21539 = 9'h9f == r_count_53_io_out ? io_r_159_b : _GEN_21538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21540 = 9'ha0 == r_count_53_io_out ? io_r_160_b : _GEN_21539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21541 = 9'ha1 == r_count_53_io_out ? io_r_161_b : _GEN_21540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21542 = 9'ha2 == r_count_53_io_out ? io_r_162_b : _GEN_21541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21543 = 9'ha3 == r_count_53_io_out ? io_r_163_b : _GEN_21542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21544 = 9'ha4 == r_count_53_io_out ? io_r_164_b : _GEN_21543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21545 = 9'ha5 == r_count_53_io_out ? io_r_165_b : _GEN_21544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21546 = 9'ha6 == r_count_53_io_out ? io_r_166_b : _GEN_21545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21547 = 9'ha7 == r_count_53_io_out ? io_r_167_b : _GEN_21546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21548 = 9'ha8 == r_count_53_io_out ? io_r_168_b : _GEN_21547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21549 = 9'ha9 == r_count_53_io_out ? io_r_169_b : _GEN_21548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21550 = 9'haa == r_count_53_io_out ? io_r_170_b : _GEN_21549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21551 = 9'hab == r_count_53_io_out ? io_r_171_b : _GEN_21550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21552 = 9'hac == r_count_53_io_out ? io_r_172_b : _GEN_21551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21553 = 9'had == r_count_53_io_out ? io_r_173_b : _GEN_21552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21554 = 9'hae == r_count_53_io_out ? io_r_174_b : _GEN_21553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21555 = 9'haf == r_count_53_io_out ? io_r_175_b : _GEN_21554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21556 = 9'hb0 == r_count_53_io_out ? io_r_176_b : _GEN_21555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21557 = 9'hb1 == r_count_53_io_out ? io_r_177_b : _GEN_21556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21558 = 9'hb2 == r_count_53_io_out ? io_r_178_b : _GEN_21557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21559 = 9'hb3 == r_count_53_io_out ? io_r_179_b : _GEN_21558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21560 = 9'hb4 == r_count_53_io_out ? io_r_180_b : _GEN_21559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21561 = 9'hb5 == r_count_53_io_out ? io_r_181_b : _GEN_21560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21562 = 9'hb6 == r_count_53_io_out ? io_r_182_b : _GEN_21561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21563 = 9'hb7 == r_count_53_io_out ? io_r_183_b : _GEN_21562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21564 = 9'hb8 == r_count_53_io_out ? io_r_184_b : _GEN_21563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21565 = 9'hb9 == r_count_53_io_out ? io_r_185_b : _GEN_21564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21566 = 9'hba == r_count_53_io_out ? io_r_186_b : _GEN_21565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21567 = 9'hbb == r_count_53_io_out ? io_r_187_b : _GEN_21566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21568 = 9'hbc == r_count_53_io_out ? io_r_188_b : _GEN_21567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21569 = 9'hbd == r_count_53_io_out ? io_r_189_b : _GEN_21568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21570 = 9'hbe == r_count_53_io_out ? io_r_190_b : _GEN_21569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21571 = 9'hbf == r_count_53_io_out ? io_r_191_b : _GEN_21570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21572 = 9'hc0 == r_count_53_io_out ? io_r_192_b : _GEN_21571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21573 = 9'hc1 == r_count_53_io_out ? io_r_193_b : _GEN_21572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21574 = 9'hc2 == r_count_53_io_out ? io_r_194_b : _GEN_21573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21575 = 9'hc3 == r_count_53_io_out ? io_r_195_b : _GEN_21574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21576 = 9'hc4 == r_count_53_io_out ? io_r_196_b : _GEN_21575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21577 = 9'hc5 == r_count_53_io_out ? io_r_197_b : _GEN_21576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21578 = 9'hc6 == r_count_53_io_out ? io_r_198_b : _GEN_21577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21579 = 9'hc7 == r_count_53_io_out ? io_r_199_b : _GEN_21578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21580 = 9'hc8 == r_count_53_io_out ? io_r_200_b : _GEN_21579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21581 = 9'hc9 == r_count_53_io_out ? io_r_201_b : _GEN_21580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21582 = 9'hca == r_count_53_io_out ? io_r_202_b : _GEN_21581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21583 = 9'hcb == r_count_53_io_out ? io_r_203_b : _GEN_21582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21584 = 9'hcc == r_count_53_io_out ? io_r_204_b : _GEN_21583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21585 = 9'hcd == r_count_53_io_out ? io_r_205_b : _GEN_21584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21586 = 9'hce == r_count_53_io_out ? io_r_206_b : _GEN_21585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21587 = 9'hcf == r_count_53_io_out ? io_r_207_b : _GEN_21586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21588 = 9'hd0 == r_count_53_io_out ? io_r_208_b : _GEN_21587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21589 = 9'hd1 == r_count_53_io_out ? io_r_209_b : _GEN_21588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21590 = 9'hd2 == r_count_53_io_out ? io_r_210_b : _GEN_21589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21591 = 9'hd3 == r_count_53_io_out ? io_r_211_b : _GEN_21590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21592 = 9'hd4 == r_count_53_io_out ? io_r_212_b : _GEN_21591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21593 = 9'hd5 == r_count_53_io_out ? io_r_213_b : _GEN_21592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21594 = 9'hd6 == r_count_53_io_out ? io_r_214_b : _GEN_21593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21595 = 9'hd7 == r_count_53_io_out ? io_r_215_b : _GEN_21594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21596 = 9'hd8 == r_count_53_io_out ? io_r_216_b : _GEN_21595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21597 = 9'hd9 == r_count_53_io_out ? io_r_217_b : _GEN_21596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21598 = 9'hda == r_count_53_io_out ? io_r_218_b : _GEN_21597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21599 = 9'hdb == r_count_53_io_out ? io_r_219_b : _GEN_21598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21600 = 9'hdc == r_count_53_io_out ? io_r_220_b : _GEN_21599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21601 = 9'hdd == r_count_53_io_out ? io_r_221_b : _GEN_21600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21602 = 9'hde == r_count_53_io_out ? io_r_222_b : _GEN_21601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21603 = 9'hdf == r_count_53_io_out ? io_r_223_b : _GEN_21602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21604 = 9'he0 == r_count_53_io_out ? io_r_224_b : _GEN_21603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21605 = 9'he1 == r_count_53_io_out ? io_r_225_b : _GEN_21604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21606 = 9'he2 == r_count_53_io_out ? io_r_226_b : _GEN_21605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21607 = 9'he3 == r_count_53_io_out ? io_r_227_b : _GEN_21606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21608 = 9'he4 == r_count_53_io_out ? io_r_228_b : _GEN_21607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21609 = 9'he5 == r_count_53_io_out ? io_r_229_b : _GEN_21608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21610 = 9'he6 == r_count_53_io_out ? io_r_230_b : _GEN_21609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21611 = 9'he7 == r_count_53_io_out ? io_r_231_b : _GEN_21610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21612 = 9'he8 == r_count_53_io_out ? io_r_232_b : _GEN_21611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21613 = 9'he9 == r_count_53_io_out ? io_r_233_b : _GEN_21612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21614 = 9'hea == r_count_53_io_out ? io_r_234_b : _GEN_21613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21615 = 9'heb == r_count_53_io_out ? io_r_235_b : _GEN_21614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21616 = 9'hec == r_count_53_io_out ? io_r_236_b : _GEN_21615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21617 = 9'hed == r_count_53_io_out ? io_r_237_b : _GEN_21616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21618 = 9'hee == r_count_53_io_out ? io_r_238_b : _GEN_21617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21619 = 9'hef == r_count_53_io_out ? io_r_239_b : _GEN_21618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21620 = 9'hf0 == r_count_53_io_out ? io_r_240_b : _GEN_21619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21621 = 9'hf1 == r_count_53_io_out ? io_r_241_b : _GEN_21620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21622 = 9'hf2 == r_count_53_io_out ? io_r_242_b : _GEN_21621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21623 = 9'hf3 == r_count_53_io_out ? io_r_243_b : _GEN_21622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21624 = 9'hf4 == r_count_53_io_out ? io_r_244_b : _GEN_21623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21625 = 9'hf5 == r_count_53_io_out ? io_r_245_b : _GEN_21624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21626 = 9'hf6 == r_count_53_io_out ? io_r_246_b : _GEN_21625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21627 = 9'hf7 == r_count_53_io_out ? io_r_247_b : _GEN_21626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21628 = 9'hf8 == r_count_53_io_out ? io_r_248_b : _GEN_21627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21629 = 9'hf9 == r_count_53_io_out ? io_r_249_b : _GEN_21628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21630 = 9'hfa == r_count_53_io_out ? io_r_250_b : _GEN_21629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21631 = 9'hfb == r_count_53_io_out ? io_r_251_b : _GEN_21630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21632 = 9'hfc == r_count_53_io_out ? io_r_252_b : _GEN_21631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21633 = 9'hfd == r_count_53_io_out ? io_r_253_b : _GEN_21632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21634 = 9'hfe == r_count_53_io_out ? io_r_254_b : _GEN_21633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21635 = 9'hff == r_count_53_io_out ? io_r_255_b : _GEN_21634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21636 = 9'h100 == r_count_53_io_out ? io_r_256_b : _GEN_21635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21637 = 9'h101 == r_count_53_io_out ? io_r_257_b : _GEN_21636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21638 = 9'h102 == r_count_53_io_out ? io_r_258_b : _GEN_21637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21639 = 9'h103 == r_count_53_io_out ? io_r_259_b : _GEN_21638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21640 = 9'h104 == r_count_53_io_out ? io_r_260_b : _GEN_21639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21641 = 9'h105 == r_count_53_io_out ? io_r_261_b : _GEN_21640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21642 = 9'h106 == r_count_53_io_out ? io_r_262_b : _GEN_21641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21643 = 9'h107 == r_count_53_io_out ? io_r_263_b : _GEN_21642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21644 = 9'h108 == r_count_53_io_out ? io_r_264_b : _GEN_21643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21645 = 9'h109 == r_count_53_io_out ? io_r_265_b : _GEN_21644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21646 = 9'h10a == r_count_53_io_out ? io_r_266_b : _GEN_21645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21647 = 9'h10b == r_count_53_io_out ? io_r_267_b : _GEN_21646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21648 = 9'h10c == r_count_53_io_out ? io_r_268_b : _GEN_21647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21649 = 9'h10d == r_count_53_io_out ? io_r_269_b : _GEN_21648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21650 = 9'h10e == r_count_53_io_out ? io_r_270_b : _GEN_21649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21651 = 9'h10f == r_count_53_io_out ? io_r_271_b : _GEN_21650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21652 = 9'h110 == r_count_53_io_out ? io_r_272_b : _GEN_21651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21653 = 9'h111 == r_count_53_io_out ? io_r_273_b : _GEN_21652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21654 = 9'h112 == r_count_53_io_out ? io_r_274_b : _GEN_21653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21655 = 9'h113 == r_count_53_io_out ? io_r_275_b : _GEN_21654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21656 = 9'h114 == r_count_53_io_out ? io_r_276_b : _GEN_21655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21657 = 9'h115 == r_count_53_io_out ? io_r_277_b : _GEN_21656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21658 = 9'h116 == r_count_53_io_out ? io_r_278_b : _GEN_21657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21659 = 9'h117 == r_count_53_io_out ? io_r_279_b : _GEN_21658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21660 = 9'h118 == r_count_53_io_out ? io_r_280_b : _GEN_21659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21661 = 9'h119 == r_count_53_io_out ? io_r_281_b : _GEN_21660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21662 = 9'h11a == r_count_53_io_out ? io_r_282_b : _GEN_21661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21663 = 9'h11b == r_count_53_io_out ? io_r_283_b : _GEN_21662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21664 = 9'h11c == r_count_53_io_out ? io_r_284_b : _GEN_21663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21665 = 9'h11d == r_count_53_io_out ? io_r_285_b : _GEN_21664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21666 = 9'h11e == r_count_53_io_out ? io_r_286_b : _GEN_21665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21667 = 9'h11f == r_count_53_io_out ? io_r_287_b : _GEN_21666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21668 = 9'h120 == r_count_53_io_out ? io_r_288_b : _GEN_21667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21669 = 9'h121 == r_count_53_io_out ? io_r_289_b : _GEN_21668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21670 = 9'h122 == r_count_53_io_out ? io_r_290_b : _GEN_21669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21671 = 9'h123 == r_count_53_io_out ? io_r_291_b : _GEN_21670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21672 = 9'h124 == r_count_53_io_out ? io_r_292_b : _GEN_21671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21673 = 9'h125 == r_count_53_io_out ? io_r_293_b : _GEN_21672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21674 = 9'h126 == r_count_53_io_out ? io_r_294_b : _GEN_21673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21675 = 9'h127 == r_count_53_io_out ? io_r_295_b : _GEN_21674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21676 = 9'h128 == r_count_53_io_out ? io_r_296_b : _GEN_21675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21677 = 9'h129 == r_count_53_io_out ? io_r_297_b : _GEN_21676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21678 = 9'h12a == r_count_53_io_out ? io_r_298_b : _GEN_21677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21679 = 9'h12b == r_count_53_io_out ? io_r_299_b : _GEN_21678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21680 = 9'h12c == r_count_53_io_out ? io_r_300_b : _GEN_21679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21681 = 9'h12d == r_count_53_io_out ? io_r_301_b : _GEN_21680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21682 = 9'h12e == r_count_53_io_out ? io_r_302_b : _GEN_21681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21683 = 9'h12f == r_count_53_io_out ? io_r_303_b : _GEN_21682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21684 = 9'h130 == r_count_53_io_out ? io_r_304_b : _GEN_21683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21685 = 9'h131 == r_count_53_io_out ? io_r_305_b : _GEN_21684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21686 = 9'h132 == r_count_53_io_out ? io_r_306_b : _GEN_21685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21687 = 9'h133 == r_count_53_io_out ? io_r_307_b : _GEN_21686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21688 = 9'h134 == r_count_53_io_out ? io_r_308_b : _GEN_21687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21689 = 9'h135 == r_count_53_io_out ? io_r_309_b : _GEN_21688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21690 = 9'h136 == r_count_53_io_out ? io_r_310_b : _GEN_21689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21691 = 9'h137 == r_count_53_io_out ? io_r_311_b : _GEN_21690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21692 = 9'h138 == r_count_53_io_out ? io_r_312_b : _GEN_21691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21693 = 9'h139 == r_count_53_io_out ? io_r_313_b : _GEN_21692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21694 = 9'h13a == r_count_53_io_out ? io_r_314_b : _GEN_21693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21695 = 9'h13b == r_count_53_io_out ? io_r_315_b : _GEN_21694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21696 = 9'h13c == r_count_53_io_out ? io_r_316_b : _GEN_21695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21697 = 9'h13d == r_count_53_io_out ? io_r_317_b : _GEN_21696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21698 = 9'h13e == r_count_53_io_out ? io_r_318_b : _GEN_21697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21699 = 9'h13f == r_count_53_io_out ? io_r_319_b : _GEN_21698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21700 = 9'h140 == r_count_53_io_out ? io_r_320_b : _GEN_21699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21701 = 9'h141 == r_count_53_io_out ? io_r_321_b : _GEN_21700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21702 = 9'h142 == r_count_53_io_out ? io_r_322_b : _GEN_21701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21703 = 9'h143 == r_count_53_io_out ? io_r_323_b : _GEN_21702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21704 = 9'h144 == r_count_53_io_out ? io_r_324_b : _GEN_21703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21705 = 9'h145 == r_count_53_io_out ? io_r_325_b : _GEN_21704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21706 = 9'h146 == r_count_53_io_out ? io_r_326_b : _GEN_21705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21707 = 9'h147 == r_count_53_io_out ? io_r_327_b : _GEN_21706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21708 = 9'h148 == r_count_53_io_out ? io_r_328_b : _GEN_21707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21709 = 9'h149 == r_count_53_io_out ? io_r_329_b : _GEN_21708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21710 = 9'h14a == r_count_53_io_out ? io_r_330_b : _GEN_21709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21711 = 9'h14b == r_count_53_io_out ? io_r_331_b : _GEN_21710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21712 = 9'h14c == r_count_53_io_out ? io_r_332_b : _GEN_21711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21713 = 9'h14d == r_count_53_io_out ? io_r_333_b : _GEN_21712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21714 = 9'h14e == r_count_53_io_out ? io_r_334_b : _GEN_21713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21715 = 9'h14f == r_count_53_io_out ? io_r_335_b : _GEN_21714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21716 = 9'h150 == r_count_53_io_out ? io_r_336_b : _GEN_21715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21717 = 9'h151 == r_count_53_io_out ? io_r_337_b : _GEN_21716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21718 = 9'h152 == r_count_53_io_out ? io_r_338_b : _GEN_21717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21719 = 9'h153 == r_count_53_io_out ? io_r_339_b : _GEN_21718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21720 = 9'h154 == r_count_53_io_out ? io_r_340_b : _GEN_21719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21721 = 9'h155 == r_count_53_io_out ? io_r_341_b : _GEN_21720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21722 = 9'h156 == r_count_53_io_out ? io_r_342_b : _GEN_21721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21723 = 9'h157 == r_count_53_io_out ? io_r_343_b : _GEN_21722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21724 = 9'h158 == r_count_53_io_out ? io_r_344_b : _GEN_21723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21725 = 9'h159 == r_count_53_io_out ? io_r_345_b : _GEN_21724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21726 = 9'h15a == r_count_53_io_out ? io_r_346_b : _GEN_21725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21727 = 9'h15b == r_count_53_io_out ? io_r_347_b : _GEN_21726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21728 = 9'h15c == r_count_53_io_out ? io_r_348_b : _GEN_21727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21729 = 9'h15d == r_count_53_io_out ? io_r_349_b : _GEN_21728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21730 = 9'h15e == r_count_53_io_out ? io_r_350_b : _GEN_21729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21731 = 9'h15f == r_count_53_io_out ? io_r_351_b : _GEN_21730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21732 = 9'h160 == r_count_53_io_out ? io_r_352_b : _GEN_21731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21733 = 9'h161 == r_count_53_io_out ? io_r_353_b : _GEN_21732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21734 = 9'h162 == r_count_53_io_out ? io_r_354_b : _GEN_21733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21735 = 9'h163 == r_count_53_io_out ? io_r_355_b : _GEN_21734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21736 = 9'h164 == r_count_53_io_out ? io_r_356_b : _GEN_21735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21737 = 9'h165 == r_count_53_io_out ? io_r_357_b : _GEN_21736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21738 = 9'h166 == r_count_53_io_out ? io_r_358_b : _GEN_21737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21739 = 9'h167 == r_count_53_io_out ? io_r_359_b : _GEN_21738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21740 = 9'h168 == r_count_53_io_out ? io_r_360_b : _GEN_21739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21741 = 9'h169 == r_count_53_io_out ? io_r_361_b : _GEN_21740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21742 = 9'h16a == r_count_53_io_out ? io_r_362_b : _GEN_21741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21743 = 9'h16b == r_count_53_io_out ? io_r_363_b : _GEN_21742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21744 = 9'h16c == r_count_53_io_out ? io_r_364_b : _GEN_21743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21745 = 9'h16d == r_count_53_io_out ? io_r_365_b : _GEN_21744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21746 = 9'h16e == r_count_53_io_out ? io_r_366_b : _GEN_21745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21747 = 9'h16f == r_count_53_io_out ? io_r_367_b : _GEN_21746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21748 = 9'h170 == r_count_53_io_out ? io_r_368_b : _GEN_21747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21749 = 9'h171 == r_count_53_io_out ? io_r_369_b : _GEN_21748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21750 = 9'h172 == r_count_53_io_out ? io_r_370_b : _GEN_21749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21751 = 9'h173 == r_count_53_io_out ? io_r_371_b : _GEN_21750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21752 = 9'h174 == r_count_53_io_out ? io_r_372_b : _GEN_21751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21753 = 9'h175 == r_count_53_io_out ? io_r_373_b : _GEN_21752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21754 = 9'h176 == r_count_53_io_out ? io_r_374_b : _GEN_21753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21755 = 9'h177 == r_count_53_io_out ? io_r_375_b : _GEN_21754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21756 = 9'h178 == r_count_53_io_out ? io_r_376_b : _GEN_21755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21757 = 9'h179 == r_count_53_io_out ? io_r_377_b : _GEN_21756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21758 = 9'h17a == r_count_53_io_out ? io_r_378_b : _GEN_21757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21759 = 9'h17b == r_count_53_io_out ? io_r_379_b : _GEN_21758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21760 = 9'h17c == r_count_53_io_out ? io_r_380_b : _GEN_21759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21761 = 9'h17d == r_count_53_io_out ? io_r_381_b : _GEN_21760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21762 = 9'h17e == r_count_53_io_out ? io_r_382_b : _GEN_21761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21763 = 9'h17f == r_count_53_io_out ? io_r_383_b : _GEN_21762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21764 = 9'h180 == r_count_53_io_out ? io_r_384_b : _GEN_21763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21765 = 9'h181 == r_count_53_io_out ? io_r_385_b : _GEN_21764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21766 = 9'h182 == r_count_53_io_out ? io_r_386_b : _GEN_21765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21767 = 9'h183 == r_count_53_io_out ? io_r_387_b : _GEN_21766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21768 = 9'h184 == r_count_53_io_out ? io_r_388_b : _GEN_21767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21769 = 9'h185 == r_count_53_io_out ? io_r_389_b : _GEN_21768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21770 = 9'h186 == r_count_53_io_out ? io_r_390_b : _GEN_21769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21771 = 9'h187 == r_count_53_io_out ? io_r_391_b : _GEN_21770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21772 = 9'h188 == r_count_53_io_out ? io_r_392_b : _GEN_21771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21773 = 9'h189 == r_count_53_io_out ? io_r_393_b : _GEN_21772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21774 = 9'h18a == r_count_53_io_out ? io_r_394_b : _GEN_21773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21775 = 9'h18b == r_count_53_io_out ? io_r_395_b : _GEN_21774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21776 = 9'h18c == r_count_53_io_out ? io_r_396_b : _GEN_21775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21777 = 9'h18d == r_count_53_io_out ? io_r_397_b : _GEN_21776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21778 = 9'h18e == r_count_53_io_out ? io_r_398_b : _GEN_21777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21781 = 9'h1 == r_count_54_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21782 = 9'h2 == r_count_54_io_out ? io_r_2_b : _GEN_21781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21783 = 9'h3 == r_count_54_io_out ? io_r_3_b : _GEN_21782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21784 = 9'h4 == r_count_54_io_out ? io_r_4_b : _GEN_21783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21785 = 9'h5 == r_count_54_io_out ? io_r_5_b : _GEN_21784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21786 = 9'h6 == r_count_54_io_out ? io_r_6_b : _GEN_21785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21787 = 9'h7 == r_count_54_io_out ? io_r_7_b : _GEN_21786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21788 = 9'h8 == r_count_54_io_out ? io_r_8_b : _GEN_21787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21789 = 9'h9 == r_count_54_io_out ? io_r_9_b : _GEN_21788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21790 = 9'ha == r_count_54_io_out ? io_r_10_b : _GEN_21789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21791 = 9'hb == r_count_54_io_out ? io_r_11_b : _GEN_21790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21792 = 9'hc == r_count_54_io_out ? io_r_12_b : _GEN_21791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21793 = 9'hd == r_count_54_io_out ? io_r_13_b : _GEN_21792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21794 = 9'he == r_count_54_io_out ? io_r_14_b : _GEN_21793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21795 = 9'hf == r_count_54_io_out ? io_r_15_b : _GEN_21794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21796 = 9'h10 == r_count_54_io_out ? io_r_16_b : _GEN_21795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21797 = 9'h11 == r_count_54_io_out ? io_r_17_b : _GEN_21796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21798 = 9'h12 == r_count_54_io_out ? io_r_18_b : _GEN_21797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21799 = 9'h13 == r_count_54_io_out ? io_r_19_b : _GEN_21798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21800 = 9'h14 == r_count_54_io_out ? io_r_20_b : _GEN_21799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21801 = 9'h15 == r_count_54_io_out ? io_r_21_b : _GEN_21800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21802 = 9'h16 == r_count_54_io_out ? io_r_22_b : _GEN_21801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21803 = 9'h17 == r_count_54_io_out ? io_r_23_b : _GEN_21802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21804 = 9'h18 == r_count_54_io_out ? io_r_24_b : _GEN_21803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21805 = 9'h19 == r_count_54_io_out ? io_r_25_b : _GEN_21804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21806 = 9'h1a == r_count_54_io_out ? io_r_26_b : _GEN_21805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21807 = 9'h1b == r_count_54_io_out ? io_r_27_b : _GEN_21806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21808 = 9'h1c == r_count_54_io_out ? io_r_28_b : _GEN_21807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21809 = 9'h1d == r_count_54_io_out ? io_r_29_b : _GEN_21808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21810 = 9'h1e == r_count_54_io_out ? io_r_30_b : _GEN_21809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21811 = 9'h1f == r_count_54_io_out ? io_r_31_b : _GEN_21810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21812 = 9'h20 == r_count_54_io_out ? io_r_32_b : _GEN_21811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21813 = 9'h21 == r_count_54_io_out ? io_r_33_b : _GEN_21812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21814 = 9'h22 == r_count_54_io_out ? io_r_34_b : _GEN_21813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21815 = 9'h23 == r_count_54_io_out ? io_r_35_b : _GEN_21814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21816 = 9'h24 == r_count_54_io_out ? io_r_36_b : _GEN_21815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21817 = 9'h25 == r_count_54_io_out ? io_r_37_b : _GEN_21816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21818 = 9'h26 == r_count_54_io_out ? io_r_38_b : _GEN_21817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21819 = 9'h27 == r_count_54_io_out ? io_r_39_b : _GEN_21818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21820 = 9'h28 == r_count_54_io_out ? io_r_40_b : _GEN_21819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21821 = 9'h29 == r_count_54_io_out ? io_r_41_b : _GEN_21820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21822 = 9'h2a == r_count_54_io_out ? io_r_42_b : _GEN_21821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21823 = 9'h2b == r_count_54_io_out ? io_r_43_b : _GEN_21822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21824 = 9'h2c == r_count_54_io_out ? io_r_44_b : _GEN_21823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21825 = 9'h2d == r_count_54_io_out ? io_r_45_b : _GEN_21824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21826 = 9'h2e == r_count_54_io_out ? io_r_46_b : _GEN_21825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21827 = 9'h2f == r_count_54_io_out ? io_r_47_b : _GEN_21826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21828 = 9'h30 == r_count_54_io_out ? io_r_48_b : _GEN_21827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21829 = 9'h31 == r_count_54_io_out ? io_r_49_b : _GEN_21828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21830 = 9'h32 == r_count_54_io_out ? io_r_50_b : _GEN_21829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21831 = 9'h33 == r_count_54_io_out ? io_r_51_b : _GEN_21830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21832 = 9'h34 == r_count_54_io_out ? io_r_52_b : _GEN_21831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21833 = 9'h35 == r_count_54_io_out ? io_r_53_b : _GEN_21832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21834 = 9'h36 == r_count_54_io_out ? io_r_54_b : _GEN_21833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21835 = 9'h37 == r_count_54_io_out ? io_r_55_b : _GEN_21834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21836 = 9'h38 == r_count_54_io_out ? io_r_56_b : _GEN_21835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21837 = 9'h39 == r_count_54_io_out ? io_r_57_b : _GEN_21836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21838 = 9'h3a == r_count_54_io_out ? io_r_58_b : _GEN_21837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21839 = 9'h3b == r_count_54_io_out ? io_r_59_b : _GEN_21838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21840 = 9'h3c == r_count_54_io_out ? io_r_60_b : _GEN_21839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21841 = 9'h3d == r_count_54_io_out ? io_r_61_b : _GEN_21840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21842 = 9'h3e == r_count_54_io_out ? io_r_62_b : _GEN_21841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21843 = 9'h3f == r_count_54_io_out ? io_r_63_b : _GEN_21842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21844 = 9'h40 == r_count_54_io_out ? io_r_64_b : _GEN_21843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21845 = 9'h41 == r_count_54_io_out ? io_r_65_b : _GEN_21844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21846 = 9'h42 == r_count_54_io_out ? io_r_66_b : _GEN_21845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21847 = 9'h43 == r_count_54_io_out ? io_r_67_b : _GEN_21846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21848 = 9'h44 == r_count_54_io_out ? io_r_68_b : _GEN_21847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21849 = 9'h45 == r_count_54_io_out ? io_r_69_b : _GEN_21848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21850 = 9'h46 == r_count_54_io_out ? io_r_70_b : _GEN_21849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21851 = 9'h47 == r_count_54_io_out ? io_r_71_b : _GEN_21850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21852 = 9'h48 == r_count_54_io_out ? io_r_72_b : _GEN_21851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21853 = 9'h49 == r_count_54_io_out ? io_r_73_b : _GEN_21852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21854 = 9'h4a == r_count_54_io_out ? io_r_74_b : _GEN_21853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21855 = 9'h4b == r_count_54_io_out ? io_r_75_b : _GEN_21854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21856 = 9'h4c == r_count_54_io_out ? io_r_76_b : _GEN_21855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21857 = 9'h4d == r_count_54_io_out ? io_r_77_b : _GEN_21856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21858 = 9'h4e == r_count_54_io_out ? io_r_78_b : _GEN_21857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21859 = 9'h4f == r_count_54_io_out ? io_r_79_b : _GEN_21858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21860 = 9'h50 == r_count_54_io_out ? io_r_80_b : _GEN_21859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21861 = 9'h51 == r_count_54_io_out ? io_r_81_b : _GEN_21860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21862 = 9'h52 == r_count_54_io_out ? io_r_82_b : _GEN_21861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21863 = 9'h53 == r_count_54_io_out ? io_r_83_b : _GEN_21862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21864 = 9'h54 == r_count_54_io_out ? io_r_84_b : _GEN_21863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21865 = 9'h55 == r_count_54_io_out ? io_r_85_b : _GEN_21864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21866 = 9'h56 == r_count_54_io_out ? io_r_86_b : _GEN_21865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21867 = 9'h57 == r_count_54_io_out ? io_r_87_b : _GEN_21866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21868 = 9'h58 == r_count_54_io_out ? io_r_88_b : _GEN_21867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21869 = 9'h59 == r_count_54_io_out ? io_r_89_b : _GEN_21868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21870 = 9'h5a == r_count_54_io_out ? io_r_90_b : _GEN_21869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21871 = 9'h5b == r_count_54_io_out ? io_r_91_b : _GEN_21870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21872 = 9'h5c == r_count_54_io_out ? io_r_92_b : _GEN_21871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21873 = 9'h5d == r_count_54_io_out ? io_r_93_b : _GEN_21872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21874 = 9'h5e == r_count_54_io_out ? io_r_94_b : _GEN_21873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21875 = 9'h5f == r_count_54_io_out ? io_r_95_b : _GEN_21874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21876 = 9'h60 == r_count_54_io_out ? io_r_96_b : _GEN_21875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21877 = 9'h61 == r_count_54_io_out ? io_r_97_b : _GEN_21876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21878 = 9'h62 == r_count_54_io_out ? io_r_98_b : _GEN_21877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21879 = 9'h63 == r_count_54_io_out ? io_r_99_b : _GEN_21878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21880 = 9'h64 == r_count_54_io_out ? io_r_100_b : _GEN_21879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21881 = 9'h65 == r_count_54_io_out ? io_r_101_b : _GEN_21880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21882 = 9'h66 == r_count_54_io_out ? io_r_102_b : _GEN_21881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21883 = 9'h67 == r_count_54_io_out ? io_r_103_b : _GEN_21882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21884 = 9'h68 == r_count_54_io_out ? io_r_104_b : _GEN_21883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21885 = 9'h69 == r_count_54_io_out ? io_r_105_b : _GEN_21884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21886 = 9'h6a == r_count_54_io_out ? io_r_106_b : _GEN_21885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21887 = 9'h6b == r_count_54_io_out ? io_r_107_b : _GEN_21886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21888 = 9'h6c == r_count_54_io_out ? io_r_108_b : _GEN_21887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21889 = 9'h6d == r_count_54_io_out ? io_r_109_b : _GEN_21888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21890 = 9'h6e == r_count_54_io_out ? io_r_110_b : _GEN_21889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21891 = 9'h6f == r_count_54_io_out ? io_r_111_b : _GEN_21890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21892 = 9'h70 == r_count_54_io_out ? io_r_112_b : _GEN_21891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21893 = 9'h71 == r_count_54_io_out ? io_r_113_b : _GEN_21892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21894 = 9'h72 == r_count_54_io_out ? io_r_114_b : _GEN_21893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21895 = 9'h73 == r_count_54_io_out ? io_r_115_b : _GEN_21894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21896 = 9'h74 == r_count_54_io_out ? io_r_116_b : _GEN_21895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21897 = 9'h75 == r_count_54_io_out ? io_r_117_b : _GEN_21896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21898 = 9'h76 == r_count_54_io_out ? io_r_118_b : _GEN_21897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21899 = 9'h77 == r_count_54_io_out ? io_r_119_b : _GEN_21898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21900 = 9'h78 == r_count_54_io_out ? io_r_120_b : _GEN_21899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21901 = 9'h79 == r_count_54_io_out ? io_r_121_b : _GEN_21900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21902 = 9'h7a == r_count_54_io_out ? io_r_122_b : _GEN_21901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21903 = 9'h7b == r_count_54_io_out ? io_r_123_b : _GEN_21902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21904 = 9'h7c == r_count_54_io_out ? io_r_124_b : _GEN_21903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21905 = 9'h7d == r_count_54_io_out ? io_r_125_b : _GEN_21904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21906 = 9'h7e == r_count_54_io_out ? io_r_126_b : _GEN_21905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21907 = 9'h7f == r_count_54_io_out ? io_r_127_b : _GEN_21906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21908 = 9'h80 == r_count_54_io_out ? io_r_128_b : _GEN_21907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21909 = 9'h81 == r_count_54_io_out ? io_r_129_b : _GEN_21908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21910 = 9'h82 == r_count_54_io_out ? io_r_130_b : _GEN_21909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21911 = 9'h83 == r_count_54_io_out ? io_r_131_b : _GEN_21910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21912 = 9'h84 == r_count_54_io_out ? io_r_132_b : _GEN_21911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21913 = 9'h85 == r_count_54_io_out ? io_r_133_b : _GEN_21912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21914 = 9'h86 == r_count_54_io_out ? io_r_134_b : _GEN_21913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21915 = 9'h87 == r_count_54_io_out ? io_r_135_b : _GEN_21914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21916 = 9'h88 == r_count_54_io_out ? io_r_136_b : _GEN_21915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21917 = 9'h89 == r_count_54_io_out ? io_r_137_b : _GEN_21916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21918 = 9'h8a == r_count_54_io_out ? io_r_138_b : _GEN_21917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21919 = 9'h8b == r_count_54_io_out ? io_r_139_b : _GEN_21918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21920 = 9'h8c == r_count_54_io_out ? io_r_140_b : _GEN_21919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21921 = 9'h8d == r_count_54_io_out ? io_r_141_b : _GEN_21920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21922 = 9'h8e == r_count_54_io_out ? io_r_142_b : _GEN_21921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21923 = 9'h8f == r_count_54_io_out ? io_r_143_b : _GEN_21922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21924 = 9'h90 == r_count_54_io_out ? io_r_144_b : _GEN_21923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21925 = 9'h91 == r_count_54_io_out ? io_r_145_b : _GEN_21924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21926 = 9'h92 == r_count_54_io_out ? io_r_146_b : _GEN_21925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21927 = 9'h93 == r_count_54_io_out ? io_r_147_b : _GEN_21926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21928 = 9'h94 == r_count_54_io_out ? io_r_148_b : _GEN_21927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21929 = 9'h95 == r_count_54_io_out ? io_r_149_b : _GEN_21928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21930 = 9'h96 == r_count_54_io_out ? io_r_150_b : _GEN_21929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21931 = 9'h97 == r_count_54_io_out ? io_r_151_b : _GEN_21930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21932 = 9'h98 == r_count_54_io_out ? io_r_152_b : _GEN_21931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21933 = 9'h99 == r_count_54_io_out ? io_r_153_b : _GEN_21932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21934 = 9'h9a == r_count_54_io_out ? io_r_154_b : _GEN_21933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21935 = 9'h9b == r_count_54_io_out ? io_r_155_b : _GEN_21934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21936 = 9'h9c == r_count_54_io_out ? io_r_156_b : _GEN_21935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21937 = 9'h9d == r_count_54_io_out ? io_r_157_b : _GEN_21936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21938 = 9'h9e == r_count_54_io_out ? io_r_158_b : _GEN_21937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21939 = 9'h9f == r_count_54_io_out ? io_r_159_b : _GEN_21938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21940 = 9'ha0 == r_count_54_io_out ? io_r_160_b : _GEN_21939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21941 = 9'ha1 == r_count_54_io_out ? io_r_161_b : _GEN_21940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21942 = 9'ha2 == r_count_54_io_out ? io_r_162_b : _GEN_21941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21943 = 9'ha3 == r_count_54_io_out ? io_r_163_b : _GEN_21942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21944 = 9'ha4 == r_count_54_io_out ? io_r_164_b : _GEN_21943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21945 = 9'ha5 == r_count_54_io_out ? io_r_165_b : _GEN_21944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21946 = 9'ha6 == r_count_54_io_out ? io_r_166_b : _GEN_21945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21947 = 9'ha7 == r_count_54_io_out ? io_r_167_b : _GEN_21946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21948 = 9'ha8 == r_count_54_io_out ? io_r_168_b : _GEN_21947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21949 = 9'ha9 == r_count_54_io_out ? io_r_169_b : _GEN_21948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21950 = 9'haa == r_count_54_io_out ? io_r_170_b : _GEN_21949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21951 = 9'hab == r_count_54_io_out ? io_r_171_b : _GEN_21950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21952 = 9'hac == r_count_54_io_out ? io_r_172_b : _GEN_21951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21953 = 9'had == r_count_54_io_out ? io_r_173_b : _GEN_21952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21954 = 9'hae == r_count_54_io_out ? io_r_174_b : _GEN_21953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21955 = 9'haf == r_count_54_io_out ? io_r_175_b : _GEN_21954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21956 = 9'hb0 == r_count_54_io_out ? io_r_176_b : _GEN_21955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21957 = 9'hb1 == r_count_54_io_out ? io_r_177_b : _GEN_21956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21958 = 9'hb2 == r_count_54_io_out ? io_r_178_b : _GEN_21957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21959 = 9'hb3 == r_count_54_io_out ? io_r_179_b : _GEN_21958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21960 = 9'hb4 == r_count_54_io_out ? io_r_180_b : _GEN_21959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21961 = 9'hb5 == r_count_54_io_out ? io_r_181_b : _GEN_21960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21962 = 9'hb6 == r_count_54_io_out ? io_r_182_b : _GEN_21961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21963 = 9'hb7 == r_count_54_io_out ? io_r_183_b : _GEN_21962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21964 = 9'hb8 == r_count_54_io_out ? io_r_184_b : _GEN_21963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21965 = 9'hb9 == r_count_54_io_out ? io_r_185_b : _GEN_21964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21966 = 9'hba == r_count_54_io_out ? io_r_186_b : _GEN_21965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21967 = 9'hbb == r_count_54_io_out ? io_r_187_b : _GEN_21966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21968 = 9'hbc == r_count_54_io_out ? io_r_188_b : _GEN_21967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21969 = 9'hbd == r_count_54_io_out ? io_r_189_b : _GEN_21968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21970 = 9'hbe == r_count_54_io_out ? io_r_190_b : _GEN_21969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21971 = 9'hbf == r_count_54_io_out ? io_r_191_b : _GEN_21970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21972 = 9'hc0 == r_count_54_io_out ? io_r_192_b : _GEN_21971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21973 = 9'hc1 == r_count_54_io_out ? io_r_193_b : _GEN_21972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21974 = 9'hc2 == r_count_54_io_out ? io_r_194_b : _GEN_21973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21975 = 9'hc3 == r_count_54_io_out ? io_r_195_b : _GEN_21974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21976 = 9'hc4 == r_count_54_io_out ? io_r_196_b : _GEN_21975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21977 = 9'hc5 == r_count_54_io_out ? io_r_197_b : _GEN_21976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21978 = 9'hc6 == r_count_54_io_out ? io_r_198_b : _GEN_21977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21979 = 9'hc7 == r_count_54_io_out ? io_r_199_b : _GEN_21978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21980 = 9'hc8 == r_count_54_io_out ? io_r_200_b : _GEN_21979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21981 = 9'hc9 == r_count_54_io_out ? io_r_201_b : _GEN_21980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21982 = 9'hca == r_count_54_io_out ? io_r_202_b : _GEN_21981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21983 = 9'hcb == r_count_54_io_out ? io_r_203_b : _GEN_21982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21984 = 9'hcc == r_count_54_io_out ? io_r_204_b : _GEN_21983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21985 = 9'hcd == r_count_54_io_out ? io_r_205_b : _GEN_21984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21986 = 9'hce == r_count_54_io_out ? io_r_206_b : _GEN_21985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21987 = 9'hcf == r_count_54_io_out ? io_r_207_b : _GEN_21986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21988 = 9'hd0 == r_count_54_io_out ? io_r_208_b : _GEN_21987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21989 = 9'hd1 == r_count_54_io_out ? io_r_209_b : _GEN_21988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21990 = 9'hd2 == r_count_54_io_out ? io_r_210_b : _GEN_21989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21991 = 9'hd3 == r_count_54_io_out ? io_r_211_b : _GEN_21990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21992 = 9'hd4 == r_count_54_io_out ? io_r_212_b : _GEN_21991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21993 = 9'hd5 == r_count_54_io_out ? io_r_213_b : _GEN_21992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21994 = 9'hd6 == r_count_54_io_out ? io_r_214_b : _GEN_21993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21995 = 9'hd7 == r_count_54_io_out ? io_r_215_b : _GEN_21994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21996 = 9'hd8 == r_count_54_io_out ? io_r_216_b : _GEN_21995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21997 = 9'hd9 == r_count_54_io_out ? io_r_217_b : _GEN_21996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21998 = 9'hda == r_count_54_io_out ? io_r_218_b : _GEN_21997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21999 = 9'hdb == r_count_54_io_out ? io_r_219_b : _GEN_21998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22000 = 9'hdc == r_count_54_io_out ? io_r_220_b : _GEN_21999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22001 = 9'hdd == r_count_54_io_out ? io_r_221_b : _GEN_22000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22002 = 9'hde == r_count_54_io_out ? io_r_222_b : _GEN_22001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22003 = 9'hdf == r_count_54_io_out ? io_r_223_b : _GEN_22002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22004 = 9'he0 == r_count_54_io_out ? io_r_224_b : _GEN_22003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22005 = 9'he1 == r_count_54_io_out ? io_r_225_b : _GEN_22004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22006 = 9'he2 == r_count_54_io_out ? io_r_226_b : _GEN_22005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22007 = 9'he3 == r_count_54_io_out ? io_r_227_b : _GEN_22006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22008 = 9'he4 == r_count_54_io_out ? io_r_228_b : _GEN_22007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22009 = 9'he5 == r_count_54_io_out ? io_r_229_b : _GEN_22008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22010 = 9'he6 == r_count_54_io_out ? io_r_230_b : _GEN_22009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22011 = 9'he7 == r_count_54_io_out ? io_r_231_b : _GEN_22010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22012 = 9'he8 == r_count_54_io_out ? io_r_232_b : _GEN_22011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22013 = 9'he9 == r_count_54_io_out ? io_r_233_b : _GEN_22012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22014 = 9'hea == r_count_54_io_out ? io_r_234_b : _GEN_22013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22015 = 9'heb == r_count_54_io_out ? io_r_235_b : _GEN_22014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22016 = 9'hec == r_count_54_io_out ? io_r_236_b : _GEN_22015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22017 = 9'hed == r_count_54_io_out ? io_r_237_b : _GEN_22016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22018 = 9'hee == r_count_54_io_out ? io_r_238_b : _GEN_22017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22019 = 9'hef == r_count_54_io_out ? io_r_239_b : _GEN_22018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22020 = 9'hf0 == r_count_54_io_out ? io_r_240_b : _GEN_22019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22021 = 9'hf1 == r_count_54_io_out ? io_r_241_b : _GEN_22020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22022 = 9'hf2 == r_count_54_io_out ? io_r_242_b : _GEN_22021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22023 = 9'hf3 == r_count_54_io_out ? io_r_243_b : _GEN_22022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22024 = 9'hf4 == r_count_54_io_out ? io_r_244_b : _GEN_22023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22025 = 9'hf5 == r_count_54_io_out ? io_r_245_b : _GEN_22024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22026 = 9'hf6 == r_count_54_io_out ? io_r_246_b : _GEN_22025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22027 = 9'hf7 == r_count_54_io_out ? io_r_247_b : _GEN_22026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22028 = 9'hf8 == r_count_54_io_out ? io_r_248_b : _GEN_22027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22029 = 9'hf9 == r_count_54_io_out ? io_r_249_b : _GEN_22028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22030 = 9'hfa == r_count_54_io_out ? io_r_250_b : _GEN_22029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22031 = 9'hfb == r_count_54_io_out ? io_r_251_b : _GEN_22030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22032 = 9'hfc == r_count_54_io_out ? io_r_252_b : _GEN_22031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22033 = 9'hfd == r_count_54_io_out ? io_r_253_b : _GEN_22032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22034 = 9'hfe == r_count_54_io_out ? io_r_254_b : _GEN_22033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22035 = 9'hff == r_count_54_io_out ? io_r_255_b : _GEN_22034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22036 = 9'h100 == r_count_54_io_out ? io_r_256_b : _GEN_22035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22037 = 9'h101 == r_count_54_io_out ? io_r_257_b : _GEN_22036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22038 = 9'h102 == r_count_54_io_out ? io_r_258_b : _GEN_22037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22039 = 9'h103 == r_count_54_io_out ? io_r_259_b : _GEN_22038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22040 = 9'h104 == r_count_54_io_out ? io_r_260_b : _GEN_22039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22041 = 9'h105 == r_count_54_io_out ? io_r_261_b : _GEN_22040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22042 = 9'h106 == r_count_54_io_out ? io_r_262_b : _GEN_22041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22043 = 9'h107 == r_count_54_io_out ? io_r_263_b : _GEN_22042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22044 = 9'h108 == r_count_54_io_out ? io_r_264_b : _GEN_22043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22045 = 9'h109 == r_count_54_io_out ? io_r_265_b : _GEN_22044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22046 = 9'h10a == r_count_54_io_out ? io_r_266_b : _GEN_22045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22047 = 9'h10b == r_count_54_io_out ? io_r_267_b : _GEN_22046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22048 = 9'h10c == r_count_54_io_out ? io_r_268_b : _GEN_22047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22049 = 9'h10d == r_count_54_io_out ? io_r_269_b : _GEN_22048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22050 = 9'h10e == r_count_54_io_out ? io_r_270_b : _GEN_22049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22051 = 9'h10f == r_count_54_io_out ? io_r_271_b : _GEN_22050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22052 = 9'h110 == r_count_54_io_out ? io_r_272_b : _GEN_22051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22053 = 9'h111 == r_count_54_io_out ? io_r_273_b : _GEN_22052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22054 = 9'h112 == r_count_54_io_out ? io_r_274_b : _GEN_22053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22055 = 9'h113 == r_count_54_io_out ? io_r_275_b : _GEN_22054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22056 = 9'h114 == r_count_54_io_out ? io_r_276_b : _GEN_22055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22057 = 9'h115 == r_count_54_io_out ? io_r_277_b : _GEN_22056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22058 = 9'h116 == r_count_54_io_out ? io_r_278_b : _GEN_22057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22059 = 9'h117 == r_count_54_io_out ? io_r_279_b : _GEN_22058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22060 = 9'h118 == r_count_54_io_out ? io_r_280_b : _GEN_22059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22061 = 9'h119 == r_count_54_io_out ? io_r_281_b : _GEN_22060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22062 = 9'h11a == r_count_54_io_out ? io_r_282_b : _GEN_22061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22063 = 9'h11b == r_count_54_io_out ? io_r_283_b : _GEN_22062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22064 = 9'h11c == r_count_54_io_out ? io_r_284_b : _GEN_22063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22065 = 9'h11d == r_count_54_io_out ? io_r_285_b : _GEN_22064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22066 = 9'h11e == r_count_54_io_out ? io_r_286_b : _GEN_22065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22067 = 9'h11f == r_count_54_io_out ? io_r_287_b : _GEN_22066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22068 = 9'h120 == r_count_54_io_out ? io_r_288_b : _GEN_22067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22069 = 9'h121 == r_count_54_io_out ? io_r_289_b : _GEN_22068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22070 = 9'h122 == r_count_54_io_out ? io_r_290_b : _GEN_22069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22071 = 9'h123 == r_count_54_io_out ? io_r_291_b : _GEN_22070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22072 = 9'h124 == r_count_54_io_out ? io_r_292_b : _GEN_22071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22073 = 9'h125 == r_count_54_io_out ? io_r_293_b : _GEN_22072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22074 = 9'h126 == r_count_54_io_out ? io_r_294_b : _GEN_22073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22075 = 9'h127 == r_count_54_io_out ? io_r_295_b : _GEN_22074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22076 = 9'h128 == r_count_54_io_out ? io_r_296_b : _GEN_22075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22077 = 9'h129 == r_count_54_io_out ? io_r_297_b : _GEN_22076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22078 = 9'h12a == r_count_54_io_out ? io_r_298_b : _GEN_22077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22079 = 9'h12b == r_count_54_io_out ? io_r_299_b : _GEN_22078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22080 = 9'h12c == r_count_54_io_out ? io_r_300_b : _GEN_22079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22081 = 9'h12d == r_count_54_io_out ? io_r_301_b : _GEN_22080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22082 = 9'h12e == r_count_54_io_out ? io_r_302_b : _GEN_22081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22083 = 9'h12f == r_count_54_io_out ? io_r_303_b : _GEN_22082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22084 = 9'h130 == r_count_54_io_out ? io_r_304_b : _GEN_22083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22085 = 9'h131 == r_count_54_io_out ? io_r_305_b : _GEN_22084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22086 = 9'h132 == r_count_54_io_out ? io_r_306_b : _GEN_22085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22087 = 9'h133 == r_count_54_io_out ? io_r_307_b : _GEN_22086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22088 = 9'h134 == r_count_54_io_out ? io_r_308_b : _GEN_22087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22089 = 9'h135 == r_count_54_io_out ? io_r_309_b : _GEN_22088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22090 = 9'h136 == r_count_54_io_out ? io_r_310_b : _GEN_22089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22091 = 9'h137 == r_count_54_io_out ? io_r_311_b : _GEN_22090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22092 = 9'h138 == r_count_54_io_out ? io_r_312_b : _GEN_22091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22093 = 9'h139 == r_count_54_io_out ? io_r_313_b : _GEN_22092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22094 = 9'h13a == r_count_54_io_out ? io_r_314_b : _GEN_22093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22095 = 9'h13b == r_count_54_io_out ? io_r_315_b : _GEN_22094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22096 = 9'h13c == r_count_54_io_out ? io_r_316_b : _GEN_22095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22097 = 9'h13d == r_count_54_io_out ? io_r_317_b : _GEN_22096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22098 = 9'h13e == r_count_54_io_out ? io_r_318_b : _GEN_22097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22099 = 9'h13f == r_count_54_io_out ? io_r_319_b : _GEN_22098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22100 = 9'h140 == r_count_54_io_out ? io_r_320_b : _GEN_22099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22101 = 9'h141 == r_count_54_io_out ? io_r_321_b : _GEN_22100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22102 = 9'h142 == r_count_54_io_out ? io_r_322_b : _GEN_22101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22103 = 9'h143 == r_count_54_io_out ? io_r_323_b : _GEN_22102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22104 = 9'h144 == r_count_54_io_out ? io_r_324_b : _GEN_22103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22105 = 9'h145 == r_count_54_io_out ? io_r_325_b : _GEN_22104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22106 = 9'h146 == r_count_54_io_out ? io_r_326_b : _GEN_22105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22107 = 9'h147 == r_count_54_io_out ? io_r_327_b : _GEN_22106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22108 = 9'h148 == r_count_54_io_out ? io_r_328_b : _GEN_22107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22109 = 9'h149 == r_count_54_io_out ? io_r_329_b : _GEN_22108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22110 = 9'h14a == r_count_54_io_out ? io_r_330_b : _GEN_22109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22111 = 9'h14b == r_count_54_io_out ? io_r_331_b : _GEN_22110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22112 = 9'h14c == r_count_54_io_out ? io_r_332_b : _GEN_22111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22113 = 9'h14d == r_count_54_io_out ? io_r_333_b : _GEN_22112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22114 = 9'h14e == r_count_54_io_out ? io_r_334_b : _GEN_22113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22115 = 9'h14f == r_count_54_io_out ? io_r_335_b : _GEN_22114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22116 = 9'h150 == r_count_54_io_out ? io_r_336_b : _GEN_22115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22117 = 9'h151 == r_count_54_io_out ? io_r_337_b : _GEN_22116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22118 = 9'h152 == r_count_54_io_out ? io_r_338_b : _GEN_22117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22119 = 9'h153 == r_count_54_io_out ? io_r_339_b : _GEN_22118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22120 = 9'h154 == r_count_54_io_out ? io_r_340_b : _GEN_22119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22121 = 9'h155 == r_count_54_io_out ? io_r_341_b : _GEN_22120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22122 = 9'h156 == r_count_54_io_out ? io_r_342_b : _GEN_22121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22123 = 9'h157 == r_count_54_io_out ? io_r_343_b : _GEN_22122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22124 = 9'h158 == r_count_54_io_out ? io_r_344_b : _GEN_22123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22125 = 9'h159 == r_count_54_io_out ? io_r_345_b : _GEN_22124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22126 = 9'h15a == r_count_54_io_out ? io_r_346_b : _GEN_22125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22127 = 9'h15b == r_count_54_io_out ? io_r_347_b : _GEN_22126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22128 = 9'h15c == r_count_54_io_out ? io_r_348_b : _GEN_22127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22129 = 9'h15d == r_count_54_io_out ? io_r_349_b : _GEN_22128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22130 = 9'h15e == r_count_54_io_out ? io_r_350_b : _GEN_22129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22131 = 9'h15f == r_count_54_io_out ? io_r_351_b : _GEN_22130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22132 = 9'h160 == r_count_54_io_out ? io_r_352_b : _GEN_22131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22133 = 9'h161 == r_count_54_io_out ? io_r_353_b : _GEN_22132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22134 = 9'h162 == r_count_54_io_out ? io_r_354_b : _GEN_22133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22135 = 9'h163 == r_count_54_io_out ? io_r_355_b : _GEN_22134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22136 = 9'h164 == r_count_54_io_out ? io_r_356_b : _GEN_22135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22137 = 9'h165 == r_count_54_io_out ? io_r_357_b : _GEN_22136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22138 = 9'h166 == r_count_54_io_out ? io_r_358_b : _GEN_22137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22139 = 9'h167 == r_count_54_io_out ? io_r_359_b : _GEN_22138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22140 = 9'h168 == r_count_54_io_out ? io_r_360_b : _GEN_22139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22141 = 9'h169 == r_count_54_io_out ? io_r_361_b : _GEN_22140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22142 = 9'h16a == r_count_54_io_out ? io_r_362_b : _GEN_22141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22143 = 9'h16b == r_count_54_io_out ? io_r_363_b : _GEN_22142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22144 = 9'h16c == r_count_54_io_out ? io_r_364_b : _GEN_22143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22145 = 9'h16d == r_count_54_io_out ? io_r_365_b : _GEN_22144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22146 = 9'h16e == r_count_54_io_out ? io_r_366_b : _GEN_22145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22147 = 9'h16f == r_count_54_io_out ? io_r_367_b : _GEN_22146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22148 = 9'h170 == r_count_54_io_out ? io_r_368_b : _GEN_22147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22149 = 9'h171 == r_count_54_io_out ? io_r_369_b : _GEN_22148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22150 = 9'h172 == r_count_54_io_out ? io_r_370_b : _GEN_22149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22151 = 9'h173 == r_count_54_io_out ? io_r_371_b : _GEN_22150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22152 = 9'h174 == r_count_54_io_out ? io_r_372_b : _GEN_22151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22153 = 9'h175 == r_count_54_io_out ? io_r_373_b : _GEN_22152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22154 = 9'h176 == r_count_54_io_out ? io_r_374_b : _GEN_22153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22155 = 9'h177 == r_count_54_io_out ? io_r_375_b : _GEN_22154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22156 = 9'h178 == r_count_54_io_out ? io_r_376_b : _GEN_22155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22157 = 9'h179 == r_count_54_io_out ? io_r_377_b : _GEN_22156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22158 = 9'h17a == r_count_54_io_out ? io_r_378_b : _GEN_22157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22159 = 9'h17b == r_count_54_io_out ? io_r_379_b : _GEN_22158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22160 = 9'h17c == r_count_54_io_out ? io_r_380_b : _GEN_22159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22161 = 9'h17d == r_count_54_io_out ? io_r_381_b : _GEN_22160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22162 = 9'h17e == r_count_54_io_out ? io_r_382_b : _GEN_22161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22163 = 9'h17f == r_count_54_io_out ? io_r_383_b : _GEN_22162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22164 = 9'h180 == r_count_54_io_out ? io_r_384_b : _GEN_22163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22165 = 9'h181 == r_count_54_io_out ? io_r_385_b : _GEN_22164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22166 = 9'h182 == r_count_54_io_out ? io_r_386_b : _GEN_22165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22167 = 9'h183 == r_count_54_io_out ? io_r_387_b : _GEN_22166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22168 = 9'h184 == r_count_54_io_out ? io_r_388_b : _GEN_22167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22169 = 9'h185 == r_count_54_io_out ? io_r_389_b : _GEN_22168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22170 = 9'h186 == r_count_54_io_out ? io_r_390_b : _GEN_22169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22171 = 9'h187 == r_count_54_io_out ? io_r_391_b : _GEN_22170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22172 = 9'h188 == r_count_54_io_out ? io_r_392_b : _GEN_22171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22173 = 9'h189 == r_count_54_io_out ? io_r_393_b : _GEN_22172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22174 = 9'h18a == r_count_54_io_out ? io_r_394_b : _GEN_22173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22175 = 9'h18b == r_count_54_io_out ? io_r_395_b : _GEN_22174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22176 = 9'h18c == r_count_54_io_out ? io_r_396_b : _GEN_22175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22177 = 9'h18d == r_count_54_io_out ? io_r_397_b : _GEN_22176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22178 = 9'h18e == r_count_54_io_out ? io_r_398_b : _GEN_22177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22181 = 9'h1 == r_count_55_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22182 = 9'h2 == r_count_55_io_out ? io_r_2_b : _GEN_22181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22183 = 9'h3 == r_count_55_io_out ? io_r_3_b : _GEN_22182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22184 = 9'h4 == r_count_55_io_out ? io_r_4_b : _GEN_22183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22185 = 9'h5 == r_count_55_io_out ? io_r_5_b : _GEN_22184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22186 = 9'h6 == r_count_55_io_out ? io_r_6_b : _GEN_22185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22187 = 9'h7 == r_count_55_io_out ? io_r_7_b : _GEN_22186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22188 = 9'h8 == r_count_55_io_out ? io_r_8_b : _GEN_22187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22189 = 9'h9 == r_count_55_io_out ? io_r_9_b : _GEN_22188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22190 = 9'ha == r_count_55_io_out ? io_r_10_b : _GEN_22189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22191 = 9'hb == r_count_55_io_out ? io_r_11_b : _GEN_22190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22192 = 9'hc == r_count_55_io_out ? io_r_12_b : _GEN_22191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22193 = 9'hd == r_count_55_io_out ? io_r_13_b : _GEN_22192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22194 = 9'he == r_count_55_io_out ? io_r_14_b : _GEN_22193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22195 = 9'hf == r_count_55_io_out ? io_r_15_b : _GEN_22194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22196 = 9'h10 == r_count_55_io_out ? io_r_16_b : _GEN_22195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22197 = 9'h11 == r_count_55_io_out ? io_r_17_b : _GEN_22196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22198 = 9'h12 == r_count_55_io_out ? io_r_18_b : _GEN_22197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22199 = 9'h13 == r_count_55_io_out ? io_r_19_b : _GEN_22198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22200 = 9'h14 == r_count_55_io_out ? io_r_20_b : _GEN_22199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22201 = 9'h15 == r_count_55_io_out ? io_r_21_b : _GEN_22200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22202 = 9'h16 == r_count_55_io_out ? io_r_22_b : _GEN_22201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22203 = 9'h17 == r_count_55_io_out ? io_r_23_b : _GEN_22202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22204 = 9'h18 == r_count_55_io_out ? io_r_24_b : _GEN_22203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22205 = 9'h19 == r_count_55_io_out ? io_r_25_b : _GEN_22204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22206 = 9'h1a == r_count_55_io_out ? io_r_26_b : _GEN_22205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22207 = 9'h1b == r_count_55_io_out ? io_r_27_b : _GEN_22206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22208 = 9'h1c == r_count_55_io_out ? io_r_28_b : _GEN_22207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22209 = 9'h1d == r_count_55_io_out ? io_r_29_b : _GEN_22208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22210 = 9'h1e == r_count_55_io_out ? io_r_30_b : _GEN_22209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22211 = 9'h1f == r_count_55_io_out ? io_r_31_b : _GEN_22210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22212 = 9'h20 == r_count_55_io_out ? io_r_32_b : _GEN_22211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22213 = 9'h21 == r_count_55_io_out ? io_r_33_b : _GEN_22212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22214 = 9'h22 == r_count_55_io_out ? io_r_34_b : _GEN_22213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22215 = 9'h23 == r_count_55_io_out ? io_r_35_b : _GEN_22214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22216 = 9'h24 == r_count_55_io_out ? io_r_36_b : _GEN_22215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22217 = 9'h25 == r_count_55_io_out ? io_r_37_b : _GEN_22216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22218 = 9'h26 == r_count_55_io_out ? io_r_38_b : _GEN_22217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22219 = 9'h27 == r_count_55_io_out ? io_r_39_b : _GEN_22218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22220 = 9'h28 == r_count_55_io_out ? io_r_40_b : _GEN_22219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22221 = 9'h29 == r_count_55_io_out ? io_r_41_b : _GEN_22220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22222 = 9'h2a == r_count_55_io_out ? io_r_42_b : _GEN_22221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22223 = 9'h2b == r_count_55_io_out ? io_r_43_b : _GEN_22222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22224 = 9'h2c == r_count_55_io_out ? io_r_44_b : _GEN_22223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22225 = 9'h2d == r_count_55_io_out ? io_r_45_b : _GEN_22224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22226 = 9'h2e == r_count_55_io_out ? io_r_46_b : _GEN_22225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22227 = 9'h2f == r_count_55_io_out ? io_r_47_b : _GEN_22226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22228 = 9'h30 == r_count_55_io_out ? io_r_48_b : _GEN_22227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22229 = 9'h31 == r_count_55_io_out ? io_r_49_b : _GEN_22228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22230 = 9'h32 == r_count_55_io_out ? io_r_50_b : _GEN_22229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22231 = 9'h33 == r_count_55_io_out ? io_r_51_b : _GEN_22230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22232 = 9'h34 == r_count_55_io_out ? io_r_52_b : _GEN_22231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22233 = 9'h35 == r_count_55_io_out ? io_r_53_b : _GEN_22232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22234 = 9'h36 == r_count_55_io_out ? io_r_54_b : _GEN_22233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22235 = 9'h37 == r_count_55_io_out ? io_r_55_b : _GEN_22234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22236 = 9'h38 == r_count_55_io_out ? io_r_56_b : _GEN_22235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22237 = 9'h39 == r_count_55_io_out ? io_r_57_b : _GEN_22236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22238 = 9'h3a == r_count_55_io_out ? io_r_58_b : _GEN_22237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22239 = 9'h3b == r_count_55_io_out ? io_r_59_b : _GEN_22238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22240 = 9'h3c == r_count_55_io_out ? io_r_60_b : _GEN_22239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22241 = 9'h3d == r_count_55_io_out ? io_r_61_b : _GEN_22240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22242 = 9'h3e == r_count_55_io_out ? io_r_62_b : _GEN_22241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22243 = 9'h3f == r_count_55_io_out ? io_r_63_b : _GEN_22242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22244 = 9'h40 == r_count_55_io_out ? io_r_64_b : _GEN_22243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22245 = 9'h41 == r_count_55_io_out ? io_r_65_b : _GEN_22244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22246 = 9'h42 == r_count_55_io_out ? io_r_66_b : _GEN_22245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22247 = 9'h43 == r_count_55_io_out ? io_r_67_b : _GEN_22246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22248 = 9'h44 == r_count_55_io_out ? io_r_68_b : _GEN_22247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22249 = 9'h45 == r_count_55_io_out ? io_r_69_b : _GEN_22248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22250 = 9'h46 == r_count_55_io_out ? io_r_70_b : _GEN_22249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22251 = 9'h47 == r_count_55_io_out ? io_r_71_b : _GEN_22250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22252 = 9'h48 == r_count_55_io_out ? io_r_72_b : _GEN_22251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22253 = 9'h49 == r_count_55_io_out ? io_r_73_b : _GEN_22252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22254 = 9'h4a == r_count_55_io_out ? io_r_74_b : _GEN_22253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22255 = 9'h4b == r_count_55_io_out ? io_r_75_b : _GEN_22254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22256 = 9'h4c == r_count_55_io_out ? io_r_76_b : _GEN_22255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22257 = 9'h4d == r_count_55_io_out ? io_r_77_b : _GEN_22256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22258 = 9'h4e == r_count_55_io_out ? io_r_78_b : _GEN_22257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22259 = 9'h4f == r_count_55_io_out ? io_r_79_b : _GEN_22258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22260 = 9'h50 == r_count_55_io_out ? io_r_80_b : _GEN_22259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22261 = 9'h51 == r_count_55_io_out ? io_r_81_b : _GEN_22260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22262 = 9'h52 == r_count_55_io_out ? io_r_82_b : _GEN_22261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22263 = 9'h53 == r_count_55_io_out ? io_r_83_b : _GEN_22262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22264 = 9'h54 == r_count_55_io_out ? io_r_84_b : _GEN_22263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22265 = 9'h55 == r_count_55_io_out ? io_r_85_b : _GEN_22264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22266 = 9'h56 == r_count_55_io_out ? io_r_86_b : _GEN_22265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22267 = 9'h57 == r_count_55_io_out ? io_r_87_b : _GEN_22266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22268 = 9'h58 == r_count_55_io_out ? io_r_88_b : _GEN_22267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22269 = 9'h59 == r_count_55_io_out ? io_r_89_b : _GEN_22268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22270 = 9'h5a == r_count_55_io_out ? io_r_90_b : _GEN_22269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22271 = 9'h5b == r_count_55_io_out ? io_r_91_b : _GEN_22270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22272 = 9'h5c == r_count_55_io_out ? io_r_92_b : _GEN_22271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22273 = 9'h5d == r_count_55_io_out ? io_r_93_b : _GEN_22272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22274 = 9'h5e == r_count_55_io_out ? io_r_94_b : _GEN_22273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22275 = 9'h5f == r_count_55_io_out ? io_r_95_b : _GEN_22274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22276 = 9'h60 == r_count_55_io_out ? io_r_96_b : _GEN_22275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22277 = 9'h61 == r_count_55_io_out ? io_r_97_b : _GEN_22276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22278 = 9'h62 == r_count_55_io_out ? io_r_98_b : _GEN_22277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22279 = 9'h63 == r_count_55_io_out ? io_r_99_b : _GEN_22278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22280 = 9'h64 == r_count_55_io_out ? io_r_100_b : _GEN_22279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22281 = 9'h65 == r_count_55_io_out ? io_r_101_b : _GEN_22280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22282 = 9'h66 == r_count_55_io_out ? io_r_102_b : _GEN_22281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22283 = 9'h67 == r_count_55_io_out ? io_r_103_b : _GEN_22282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22284 = 9'h68 == r_count_55_io_out ? io_r_104_b : _GEN_22283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22285 = 9'h69 == r_count_55_io_out ? io_r_105_b : _GEN_22284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22286 = 9'h6a == r_count_55_io_out ? io_r_106_b : _GEN_22285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22287 = 9'h6b == r_count_55_io_out ? io_r_107_b : _GEN_22286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22288 = 9'h6c == r_count_55_io_out ? io_r_108_b : _GEN_22287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22289 = 9'h6d == r_count_55_io_out ? io_r_109_b : _GEN_22288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22290 = 9'h6e == r_count_55_io_out ? io_r_110_b : _GEN_22289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22291 = 9'h6f == r_count_55_io_out ? io_r_111_b : _GEN_22290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22292 = 9'h70 == r_count_55_io_out ? io_r_112_b : _GEN_22291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22293 = 9'h71 == r_count_55_io_out ? io_r_113_b : _GEN_22292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22294 = 9'h72 == r_count_55_io_out ? io_r_114_b : _GEN_22293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22295 = 9'h73 == r_count_55_io_out ? io_r_115_b : _GEN_22294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22296 = 9'h74 == r_count_55_io_out ? io_r_116_b : _GEN_22295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22297 = 9'h75 == r_count_55_io_out ? io_r_117_b : _GEN_22296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22298 = 9'h76 == r_count_55_io_out ? io_r_118_b : _GEN_22297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22299 = 9'h77 == r_count_55_io_out ? io_r_119_b : _GEN_22298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22300 = 9'h78 == r_count_55_io_out ? io_r_120_b : _GEN_22299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22301 = 9'h79 == r_count_55_io_out ? io_r_121_b : _GEN_22300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22302 = 9'h7a == r_count_55_io_out ? io_r_122_b : _GEN_22301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22303 = 9'h7b == r_count_55_io_out ? io_r_123_b : _GEN_22302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22304 = 9'h7c == r_count_55_io_out ? io_r_124_b : _GEN_22303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22305 = 9'h7d == r_count_55_io_out ? io_r_125_b : _GEN_22304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22306 = 9'h7e == r_count_55_io_out ? io_r_126_b : _GEN_22305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22307 = 9'h7f == r_count_55_io_out ? io_r_127_b : _GEN_22306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22308 = 9'h80 == r_count_55_io_out ? io_r_128_b : _GEN_22307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22309 = 9'h81 == r_count_55_io_out ? io_r_129_b : _GEN_22308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22310 = 9'h82 == r_count_55_io_out ? io_r_130_b : _GEN_22309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22311 = 9'h83 == r_count_55_io_out ? io_r_131_b : _GEN_22310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22312 = 9'h84 == r_count_55_io_out ? io_r_132_b : _GEN_22311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22313 = 9'h85 == r_count_55_io_out ? io_r_133_b : _GEN_22312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22314 = 9'h86 == r_count_55_io_out ? io_r_134_b : _GEN_22313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22315 = 9'h87 == r_count_55_io_out ? io_r_135_b : _GEN_22314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22316 = 9'h88 == r_count_55_io_out ? io_r_136_b : _GEN_22315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22317 = 9'h89 == r_count_55_io_out ? io_r_137_b : _GEN_22316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22318 = 9'h8a == r_count_55_io_out ? io_r_138_b : _GEN_22317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22319 = 9'h8b == r_count_55_io_out ? io_r_139_b : _GEN_22318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22320 = 9'h8c == r_count_55_io_out ? io_r_140_b : _GEN_22319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22321 = 9'h8d == r_count_55_io_out ? io_r_141_b : _GEN_22320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22322 = 9'h8e == r_count_55_io_out ? io_r_142_b : _GEN_22321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22323 = 9'h8f == r_count_55_io_out ? io_r_143_b : _GEN_22322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22324 = 9'h90 == r_count_55_io_out ? io_r_144_b : _GEN_22323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22325 = 9'h91 == r_count_55_io_out ? io_r_145_b : _GEN_22324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22326 = 9'h92 == r_count_55_io_out ? io_r_146_b : _GEN_22325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22327 = 9'h93 == r_count_55_io_out ? io_r_147_b : _GEN_22326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22328 = 9'h94 == r_count_55_io_out ? io_r_148_b : _GEN_22327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22329 = 9'h95 == r_count_55_io_out ? io_r_149_b : _GEN_22328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22330 = 9'h96 == r_count_55_io_out ? io_r_150_b : _GEN_22329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22331 = 9'h97 == r_count_55_io_out ? io_r_151_b : _GEN_22330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22332 = 9'h98 == r_count_55_io_out ? io_r_152_b : _GEN_22331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22333 = 9'h99 == r_count_55_io_out ? io_r_153_b : _GEN_22332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22334 = 9'h9a == r_count_55_io_out ? io_r_154_b : _GEN_22333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22335 = 9'h9b == r_count_55_io_out ? io_r_155_b : _GEN_22334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22336 = 9'h9c == r_count_55_io_out ? io_r_156_b : _GEN_22335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22337 = 9'h9d == r_count_55_io_out ? io_r_157_b : _GEN_22336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22338 = 9'h9e == r_count_55_io_out ? io_r_158_b : _GEN_22337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22339 = 9'h9f == r_count_55_io_out ? io_r_159_b : _GEN_22338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22340 = 9'ha0 == r_count_55_io_out ? io_r_160_b : _GEN_22339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22341 = 9'ha1 == r_count_55_io_out ? io_r_161_b : _GEN_22340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22342 = 9'ha2 == r_count_55_io_out ? io_r_162_b : _GEN_22341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22343 = 9'ha3 == r_count_55_io_out ? io_r_163_b : _GEN_22342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22344 = 9'ha4 == r_count_55_io_out ? io_r_164_b : _GEN_22343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22345 = 9'ha5 == r_count_55_io_out ? io_r_165_b : _GEN_22344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22346 = 9'ha6 == r_count_55_io_out ? io_r_166_b : _GEN_22345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22347 = 9'ha7 == r_count_55_io_out ? io_r_167_b : _GEN_22346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22348 = 9'ha8 == r_count_55_io_out ? io_r_168_b : _GEN_22347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22349 = 9'ha9 == r_count_55_io_out ? io_r_169_b : _GEN_22348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22350 = 9'haa == r_count_55_io_out ? io_r_170_b : _GEN_22349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22351 = 9'hab == r_count_55_io_out ? io_r_171_b : _GEN_22350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22352 = 9'hac == r_count_55_io_out ? io_r_172_b : _GEN_22351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22353 = 9'had == r_count_55_io_out ? io_r_173_b : _GEN_22352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22354 = 9'hae == r_count_55_io_out ? io_r_174_b : _GEN_22353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22355 = 9'haf == r_count_55_io_out ? io_r_175_b : _GEN_22354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22356 = 9'hb0 == r_count_55_io_out ? io_r_176_b : _GEN_22355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22357 = 9'hb1 == r_count_55_io_out ? io_r_177_b : _GEN_22356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22358 = 9'hb2 == r_count_55_io_out ? io_r_178_b : _GEN_22357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22359 = 9'hb3 == r_count_55_io_out ? io_r_179_b : _GEN_22358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22360 = 9'hb4 == r_count_55_io_out ? io_r_180_b : _GEN_22359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22361 = 9'hb5 == r_count_55_io_out ? io_r_181_b : _GEN_22360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22362 = 9'hb6 == r_count_55_io_out ? io_r_182_b : _GEN_22361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22363 = 9'hb7 == r_count_55_io_out ? io_r_183_b : _GEN_22362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22364 = 9'hb8 == r_count_55_io_out ? io_r_184_b : _GEN_22363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22365 = 9'hb9 == r_count_55_io_out ? io_r_185_b : _GEN_22364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22366 = 9'hba == r_count_55_io_out ? io_r_186_b : _GEN_22365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22367 = 9'hbb == r_count_55_io_out ? io_r_187_b : _GEN_22366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22368 = 9'hbc == r_count_55_io_out ? io_r_188_b : _GEN_22367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22369 = 9'hbd == r_count_55_io_out ? io_r_189_b : _GEN_22368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22370 = 9'hbe == r_count_55_io_out ? io_r_190_b : _GEN_22369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22371 = 9'hbf == r_count_55_io_out ? io_r_191_b : _GEN_22370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22372 = 9'hc0 == r_count_55_io_out ? io_r_192_b : _GEN_22371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22373 = 9'hc1 == r_count_55_io_out ? io_r_193_b : _GEN_22372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22374 = 9'hc2 == r_count_55_io_out ? io_r_194_b : _GEN_22373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22375 = 9'hc3 == r_count_55_io_out ? io_r_195_b : _GEN_22374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22376 = 9'hc4 == r_count_55_io_out ? io_r_196_b : _GEN_22375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22377 = 9'hc5 == r_count_55_io_out ? io_r_197_b : _GEN_22376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22378 = 9'hc6 == r_count_55_io_out ? io_r_198_b : _GEN_22377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22379 = 9'hc7 == r_count_55_io_out ? io_r_199_b : _GEN_22378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22380 = 9'hc8 == r_count_55_io_out ? io_r_200_b : _GEN_22379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22381 = 9'hc9 == r_count_55_io_out ? io_r_201_b : _GEN_22380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22382 = 9'hca == r_count_55_io_out ? io_r_202_b : _GEN_22381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22383 = 9'hcb == r_count_55_io_out ? io_r_203_b : _GEN_22382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22384 = 9'hcc == r_count_55_io_out ? io_r_204_b : _GEN_22383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22385 = 9'hcd == r_count_55_io_out ? io_r_205_b : _GEN_22384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22386 = 9'hce == r_count_55_io_out ? io_r_206_b : _GEN_22385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22387 = 9'hcf == r_count_55_io_out ? io_r_207_b : _GEN_22386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22388 = 9'hd0 == r_count_55_io_out ? io_r_208_b : _GEN_22387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22389 = 9'hd1 == r_count_55_io_out ? io_r_209_b : _GEN_22388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22390 = 9'hd2 == r_count_55_io_out ? io_r_210_b : _GEN_22389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22391 = 9'hd3 == r_count_55_io_out ? io_r_211_b : _GEN_22390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22392 = 9'hd4 == r_count_55_io_out ? io_r_212_b : _GEN_22391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22393 = 9'hd5 == r_count_55_io_out ? io_r_213_b : _GEN_22392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22394 = 9'hd6 == r_count_55_io_out ? io_r_214_b : _GEN_22393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22395 = 9'hd7 == r_count_55_io_out ? io_r_215_b : _GEN_22394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22396 = 9'hd8 == r_count_55_io_out ? io_r_216_b : _GEN_22395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22397 = 9'hd9 == r_count_55_io_out ? io_r_217_b : _GEN_22396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22398 = 9'hda == r_count_55_io_out ? io_r_218_b : _GEN_22397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22399 = 9'hdb == r_count_55_io_out ? io_r_219_b : _GEN_22398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22400 = 9'hdc == r_count_55_io_out ? io_r_220_b : _GEN_22399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22401 = 9'hdd == r_count_55_io_out ? io_r_221_b : _GEN_22400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22402 = 9'hde == r_count_55_io_out ? io_r_222_b : _GEN_22401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22403 = 9'hdf == r_count_55_io_out ? io_r_223_b : _GEN_22402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22404 = 9'he0 == r_count_55_io_out ? io_r_224_b : _GEN_22403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22405 = 9'he1 == r_count_55_io_out ? io_r_225_b : _GEN_22404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22406 = 9'he2 == r_count_55_io_out ? io_r_226_b : _GEN_22405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22407 = 9'he3 == r_count_55_io_out ? io_r_227_b : _GEN_22406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22408 = 9'he4 == r_count_55_io_out ? io_r_228_b : _GEN_22407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22409 = 9'he5 == r_count_55_io_out ? io_r_229_b : _GEN_22408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22410 = 9'he6 == r_count_55_io_out ? io_r_230_b : _GEN_22409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22411 = 9'he7 == r_count_55_io_out ? io_r_231_b : _GEN_22410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22412 = 9'he8 == r_count_55_io_out ? io_r_232_b : _GEN_22411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22413 = 9'he9 == r_count_55_io_out ? io_r_233_b : _GEN_22412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22414 = 9'hea == r_count_55_io_out ? io_r_234_b : _GEN_22413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22415 = 9'heb == r_count_55_io_out ? io_r_235_b : _GEN_22414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22416 = 9'hec == r_count_55_io_out ? io_r_236_b : _GEN_22415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22417 = 9'hed == r_count_55_io_out ? io_r_237_b : _GEN_22416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22418 = 9'hee == r_count_55_io_out ? io_r_238_b : _GEN_22417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22419 = 9'hef == r_count_55_io_out ? io_r_239_b : _GEN_22418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22420 = 9'hf0 == r_count_55_io_out ? io_r_240_b : _GEN_22419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22421 = 9'hf1 == r_count_55_io_out ? io_r_241_b : _GEN_22420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22422 = 9'hf2 == r_count_55_io_out ? io_r_242_b : _GEN_22421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22423 = 9'hf3 == r_count_55_io_out ? io_r_243_b : _GEN_22422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22424 = 9'hf4 == r_count_55_io_out ? io_r_244_b : _GEN_22423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22425 = 9'hf5 == r_count_55_io_out ? io_r_245_b : _GEN_22424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22426 = 9'hf6 == r_count_55_io_out ? io_r_246_b : _GEN_22425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22427 = 9'hf7 == r_count_55_io_out ? io_r_247_b : _GEN_22426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22428 = 9'hf8 == r_count_55_io_out ? io_r_248_b : _GEN_22427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22429 = 9'hf9 == r_count_55_io_out ? io_r_249_b : _GEN_22428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22430 = 9'hfa == r_count_55_io_out ? io_r_250_b : _GEN_22429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22431 = 9'hfb == r_count_55_io_out ? io_r_251_b : _GEN_22430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22432 = 9'hfc == r_count_55_io_out ? io_r_252_b : _GEN_22431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22433 = 9'hfd == r_count_55_io_out ? io_r_253_b : _GEN_22432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22434 = 9'hfe == r_count_55_io_out ? io_r_254_b : _GEN_22433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22435 = 9'hff == r_count_55_io_out ? io_r_255_b : _GEN_22434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22436 = 9'h100 == r_count_55_io_out ? io_r_256_b : _GEN_22435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22437 = 9'h101 == r_count_55_io_out ? io_r_257_b : _GEN_22436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22438 = 9'h102 == r_count_55_io_out ? io_r_258_b : _GEN_22437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22439 = 9'h103 == r_count_55_io_out ? io_r_259_b : _GEN_22438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22440 = 9'h104 == r_count_55_io_out ? io_r_260_b : _GEN_22439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22441 = 9'h105 == r_count_55_io_out ? io_r_261_b : _GEN_22440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22442 = 9'h106 == r_count_55_io_out ? io_r_262_b : _GEN_22441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22443 = 9'h107 == r_count_55_io_out ? io_r_263_b : _GEN_22442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22444 = 9'h108 == r_count_55_io_out ? io_r_264_b : _GEN_22443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22445 = 9'h109 == r_count_55_io_out ? io_r_265_b : _GEN_22444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22446 = 9'h10a == r_count_55_io_out ? io_r_266_b : _GEN_22445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22447 = 9'h10b == r_count_55_io_out ? io_r_267_b : _GEN_22446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22448 = 9'h10c == r_count_55_io_out ? io_r_268_b : _GEN_22447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22449 = 9'h10d == r_count_55_io_out ? io_r_269_b : _GEN_22448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22450 = 9'h10e == r_count_55_io_out ? io_r_270_b : _GEN_22449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22451 = 9'h10f == r_count_55_io_out ? io_r_271_b : _GEN_22450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22452 = 9'h110 == r_count_55_io_out ? io_r_272_b : _GEN_22451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22453 = 9'h111 == r_count_55_io_out ? io_r_273_b : _GEN_22452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22454 = 9'h112 == r_count_55_io_out ? io_r_274_b : _GEN_22453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22455 = 9'h113 == r_count_55_io_out ? io_r_275_b : _GEN_22454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22456 = 9'h114 == r_count_55_io_out ? io_r_276_b : _GEN_22455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22457 = 9'h115 == r_count_55_io_out ? io_r_277_b : _GEN_22456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22458 = 9'h116 == r_count_55_io_out ? io_r_278_b : _GEN_22457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22459 = 9'h117 == r_count_55_io_out ? io_r_279_b : _GEN_22458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22460 = 9'h118 == r_count_55_io_out ? io_r_280_b : _GEN_22459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22461 = 9'h119 == r_count_55_io_out ? io_r_281_b : _GEN_22460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22462 = 9'h11a == r_count_55_io_out ? io_r_282_b : _GEN_22461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22463 = 9'h11b == r_count_55_io_out ? io_r_283_b : _GEN_22462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22464 = 9'h11c == r_count_55_io_out ? io_r_284_b : _GEN_22463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22465 = 9'h11d == r_count_55_io_out ? io_r_285_b : _GEN_22464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22466 = 9'h11e == r_count_55_io_out ? io_r_286_b : _GEN_22465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22467 = 9'h11f == r_count_55_io_out ? io_r_287_b : _GEN_22466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22468 = 9'h120 == r_count_55_io_out ? io_r_288_b : _GEN_22467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22469 = 9'h121 == r_count_55_io_out ? io_r_289_b : _GEN_22468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22470 = 9'h122 == r_count_55_io_out ? io_r_290_b : _GEN_22469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22471 = 9'h123 == r_count_55_io_out ? io_r_291_b : _GEN_22470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22472 = 9'h124 == r_count_55_io_out ? io_r_292_b : _GEN_22471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22473 = 9'h125 == r_count_55_io_out ? io_r_293_b : _GEN_22472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22474 = 9'h126 == r_count_55_io_out ? io_r_294_b : _GEN_22473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22475 = 9'h127 == r_count_55_io_out ? io_r_295_b : _GEN_22474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22476 = 9'h128 == r_count_55_io_out ? io_r_296_b : _GEN_22475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22477 = 9'h129 == r_count_55_io_out ? io_r_297_b : _GEN_22476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22478 = 9'h12a == r_count_55_io_out ? io_r_298_b : _GEN_22477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22479 = 9'h12b == r_count_55_io_out ? io_r_299_b : _GEN_22478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22480 = 9'h12c == r_count_55_io_out ? io_r_300_b : _GEN_22479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22481 = 9'h12d == r_count_55_io_out ? io_r_301_b : _GEN_22480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22482 = 9'h12e == r_count_55_io_out ? io_r_302_b : _GEN_22481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22483 = 9'h12f == r_count_55_io_out ? io_r_303_b : _GEN_22482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22484 = 9'h130 == r_count_55_io_out ? io_r_304_b : _GEN_22483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22485 = 9'h131 == r_count_55_io_out ? io_r_305_b : _GEN_22484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22486 = 9'h132 == r_count_55_io_out ? io_r_306_b : _GEN_22485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22487 = 9'h133 == r_count_55_io_out ? io_r_307_b : _GEN_22486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22488 = 9'h134 == r_count_55_io_out ? io_r_308_b : _GEN_22487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22489 = 9'h135 == r_count_55_io_out ? io_r_309_b : _GEN_22488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22490 = 9'h136 == r_count_55_io_out ? io_r_310_b : _GEN_22489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22491 = 9'h137 == r_count_55_io_out ? io_r_311_b : _GEN_22490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22492 = 9'h138 == r_count_55_io_out ? io_r_312_b : _GEN_22491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22493 = 9'h139 == r_count_55_io_out ? io_r_313_b : _GEN_22492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22494 = 9'h13a == r_count_55_io_out ? io_r_314_b : _GEN_22493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22495 = 9'h13b == r_count_55_io_out ? io_r_315_b : _GEN_22494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22496 = 9'h13c == r_count_55_io_out ? io_r_316_b : _GEN_22495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22497 = 9'h13d == r_count_55_io_out ? io_r_317_b : _GEN_22496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22498 = 9'h13e == r_count_55_io_out ? io_r_318_b : _GEN_22497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22499 = 9'h13f == r_count_55_io_out ? io_r_319_b : _GEN_22498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22500 = 9'h140 == r_count_55_io_out ? io_r_320_b : _GEN_22499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22501 = 9'h141 == r_count_55_io_out ? io_r_321_b : _GEN_22500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22502 = 9'h142 == r_count_55_io_out ? io_r_322_b : _GEN_22501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22503 = 9'h143 == r_count_55_io_out ? io_r_323_b : _GEN_22502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22504 = 9'h144 == r_count_55_io_out ? io_r_324_b : _GEN_22503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22505 = 9'h145 == r_count_55_io_out ? io_r_325_b : _GEN_22504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22506 = 9'h146 == r_count_55_io_out ? io_r_326_b : _GEN_22505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22507 = 9'h147 == r_count_55_io_out ? io_r_327_b : _GEN_22506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22508 = 9'h148 == r_count_55_io_out ? io_r_328_b : _GEN_22507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22509 = 9'h149 == r_count_55_io_out ? io_r_329_b : _GEN_22508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22510 = 9'h14a == r_count_55_io_out ? io_r_330_b : _GEN_22509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22511 = 9'h14b == r_count_55_io_out ? io_r_331_b : _GEN_22510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22512 = 9'h14c == r_count_55_io_out ? io_r_332_b : _GEN_22511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22513 = 9'h14d == r_count_55_io_out ? io_r_333_b : _GEN_22512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22514 = 9'h14e == r_count_55_io_out ? io_r_334_b : _GEN_22513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22515 = 9'h14f == r_count_55_io_out ? io_r_335_b : _GEN_22514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22516 = 9'h150 == r_count_55_io_out ? io_r_336_b : _GEN_22515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22517 = 9'h151 == r_count_55_io_out ? io_r_337_b : _GEN_22516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22518 = 9'h152 == r_count_55_io_out ? io_r_338_b : _GEN_22517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22519 = 9'h153 == r_count_55_io_out ? io_r_339_b : _GEN_22518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22520 = 9'h154 == r_count_55_io_out ? io_r_340_b : _GEN_22519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22521 = 9'h155 == r_count_55_io_out ? io_r_341_b : _GEN_22520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22522 = 9'h156 == r_count_55_io_out ? io_r_342_b : _GEN_22521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22523 = 9'h157 == r_count_55_io_out ? io_r_343_b : _GEN_22522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22524 = 9'h158 == r_count_55_io_out ? io_r_344_b : _GEN_22523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22525 = 9'h159 == r_count_55_io_out ? io_r_345_b : _GEN_22524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22526 = 9'h15a == r_count_55_io_out ? io_r_346_b : _GEN_22525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22527 = 9'h15b == r_count_55_io_out ? io_r_347_b : _GEN_22526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22528 = 9'h15c == r_count_55_io_out ? io_r_348_b : _GEN_22527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22529 = 9'h15d == r_count_55_io_out ? io_r_349_b : _GEN_22528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22530 = 9'h15e == r_count_55_io_out ? io_r_350_b : _GEN_22529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22531 = 9'h15f == r_count_55_io_out ? io_r_351_b : _GEN_22530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22532 = 9'h160 == r_count_55_io_out ? io_r_352_b : _GEN_22531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22533 = 9'h161 == r_count_55_io_out ? io_r_353_b : _GEN_22532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22534 = 9'h162 == r_count_55_io_out ? io_r_354_b : _GEN_22533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22535 = 9'h163 == r_count_55_io_out ? io_r_355_b : _GEN_22534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22536 = 9'h164 == r_count_55_io_out ? io_r_356_b : _GEN_22535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22537 = 9'h165 == r_count_55_io_out ? io_r_357_b : _GEN_22536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22538 = 9'h166 == r_count_55_io_out ? io_r_358_b : _GEN_22537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22539 = 9'h167 == r_count_55_io_out ? io_r_359_b : _GEN_22538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22540 = 9'h168 == r_count_55_io_out ? io_r_360_b : _GEN_22539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22541 = 9'h169 == r_count_55_io_out ? io_r_361_b : _GEN_22540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22542 = 9'h16a == r_count_55_io_out ? io_r_362_b : _GEN_22541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22543 = 9'h16b == r_count_55_io_out ? io_r_363_b : _GEN_22542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22544 = 9'h16c == r_count_55_io_out ? io_r_364_b : _GEN_22543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22545 = 9'h16d == r_count_55_io_out ? io_r_365_b : _GEN_22544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22546 = 9'h16e == r_count_55_io_out ? io_r_366_b : _GEN_22545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22547 = 9'h16f == r_count_55_io_out ? io_r_367_b : _GEN_22546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22548 = 9'h170 == r_count_55_io_out ? io_r_368_b : _GEN_22547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22549 = 9'h171 == r_count_55_io_out ? io_r_369_b : _GEN_22548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22550 = 9'h172 == r_count_55_io_out ? io_r_370_b : _GEN_22549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22551 = 9'h173 == r_count_55_io_out ? io_r_371_b : _GEN_22550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22552 = 9'h174 == r_count_55_io_out ? io_r_372_b : _GEN_22551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22553 = 9'h175 == r_count_55_io_out ? io_r_373_b : _GEN_22552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22554 = 9'h176 == r_count_55_io_out ? io_r_374_b : _GEN_22553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22555 = 9'h177 == r_count_55_io_out ? io_r_375_b : _GEN_22554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22556 = 9'h178 == r_count_55_io_out ? io_r_376_b : _GEN_22555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22557 = 9'h179 == r_count_55_io_out ? io_r_377_b : _GEN_22556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22558 = 9'h17a == r_count_55_io_out ? io_r_378_b : _GEN_22557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22559 = 9'h17b == r_count_55_io_out ? io_r_379_b : _GEN_22558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22560 = 9'h17c == r_count_55_io_out ? io_r_380_b : _GEN_22559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22561 = 9'h17d == r_count_55_io_out ? io_r_381_b : _GEN_22560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22562 = 9'h17e == r_count_55_io_out ? io_r_382_b : _GEN_22561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22563 = 9'h17f == r_count_55_io_out ? io_r_383_b : _GEN_22562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22564 = 9'h180 == r_count_55_io_out ? io_r_384_b : _GEN_22563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22565 = 9'h181 == r_count_55_io_out ? io_r_385_b : _GEN_22564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22566 = 9'h182 == r_count_55_io_out ? io_r_386_b : _GEN_22565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22567 = 9'h183 == r_count_55_io_out ? io_r_387_b : _GEN_22566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22568 = 9'h184 == r_count_55_io_out ? io_r_388_b : _GEN_22567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22569 = 9'h185 == r_count_55_io_out ? io_r_389_b : _GEN_22568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22570 = 9'h186 == r_count_55_io_out ? io_r_390_b : _GEN_22569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22571 = 9'h187 == r_count_55_io_out ? io_r_391_b : _GEN_22570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22572 = 9'h188 == r_count_55_io_out ? io_r_392_b : _GEN_22571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22573 = 9'h189 == r_count_55_io_out ? io_r_393_b : _GEN_22572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22574 = 9'h18a == r_count_55_io_out ? io_r_394_b : _GEN_22573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22575 = 9'h18b == r_count_55_io_out ? io_r_395_b : _GEN_22574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22576 = 9'h18c == r_count_55_io_out ? io_r_396_b : _GEN_22575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22577 = 9'h18d == r_count_55_io_out ? io_r_397_b : _GEN_22576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22578 = 9'h18e == r_count_55_io_out ? io_r_398_b : _GEN_22577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22581 = 9'h1 == r_count_56_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22582 = 9'h2 == r_count_56_io_out ? io_r_2_b : _GEN_22581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22583 = 9'h3 == r_count_56_io_out ? io_r_3_b : _GEN_22582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22584 = 9'h4 == r_count_56_io_out ? io_r_4_b : _GEN_22583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22585 = 9'h5 == r_count_56_io_out ? io_r_5_b : _GEN_22584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22586 = 9'h6 == r_count_56_io_out ? io_r_6_b : _GEN_22585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22587 = 9'h7 == r_count_56_io_out ? io_r_7_b : _GEN_22586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22588 = 9'h8 == r_count_56_io_out ? io_r_8_b : _GEN_22587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22589 = 9'h9 == r_count_56_io_out ? io_r_9_b : _GEN_22588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22590 = 9'ha == r_count_56_io_out ? io_r_10_b : _GEN_22589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22591 = 9'hb == r_count_56_io_out ? io_r_11_b : _GEN_22590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22592 = 9'hc == r_count_56_io_out ? io_r_12_b : _GEN_22591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22593 = 9'hd == r_count_56_io_out ? io_r_13_b : _GEN_22592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22594 = 9'he == r_count_56_io_out ? io_r_14_b : _GEN_22593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22595 = 9'hf == r_count_56_io_out ? io_r_15_b : _GEN_22594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22596 = 9'h10 == r_count_56_io_out ? io_r_16_b : _GEN_22595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22597 = 9'h11 == r_count_56_io_out ? io_r_17_b : _GEN_22596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22598 = 9'h12 == r_count_56_io_out ? io_r_18_b : _GEN_22597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22599 = 9'h13 == r_count_56_io_out ? io_r_19_b : _GEN_22598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22600 = 9'h14 == r_count_56_io_out ? io_r_20_b : _GEN_22599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22601 = 9'h15 == r_count_56_io_out ? io_r_21_b : _GEN_22600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22602 = 9'h16 == r_count_56_io_out ? io_r_22_b : _GEN_22601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22603 = 9'h17 == r_count_56_io_out ? io_r_23_b : _GEN_22602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22604 = 9'h18 == r_count_56_io_out ? io_r_24_b : _GEN_22603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22605 = 9'h19 == r_count_56_io_out ? io_r_25_b : _GEN_22604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22606 = 9'h1a == r_count_56_io_out ? io_r_26_b : _GEN_22605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22607 = 9'h1b == r_count_56_io_out ? io_r_27_b : _GEN_22606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22608 = 9'h1c == r_count_56_io_out ? io_r_28_b : _GEN_22607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22609 = 9'h1d == r_count_56_io_out ? io_r_29_b : _GEN_22608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22610 = 9'h1e == r_count_56_io_out ? io_r_30_b : _GEN_22609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22611 = 9'h1f == r_count_56_io_out ? io_r_31_b : _GEN_22610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22612 = 9'h20 == r_count_56_io_out ? io_r_32_b : _GEN_22611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22613 = 9'h21 == r_count_56_io_out ? io_r_33_b : _GEN_22612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22614 = 9'h22 == r_count_56_io_out ? io_r_34_b : _GEN_22613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22615 = 9'h23 == r_count_56_io_out ? io_r_35_b : _GEN_22614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22616 = 9'h24 == r_count_56_io_out ? io_r_36_b : _GEN_22615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22617 = 9'h25 == r_count_56_io_out ? io_r_37_b : _GEN_22616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22618 = 9'h26 == r_count_56_io_out ? io_r_38_b : _GEN_22617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22619 = 9'h27 == r_count_56_io_out ? io_r_39_b : _GEN_22618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22620 = 9'h28 == r_count_56_io_out ? io_r_40_b : _GEN_22619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22621 = 9'h29 == r_count_56_io_out ? io_r_41_b : _GEN_22620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22622 = 9'h2a == r_count_56_io_out ? io_r_42_b : _GEN_22621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22623 = 9'h2b == r_count_56_io_out ? io_r_43_b : _GEN_22622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22624 = 9'h2c == r_count_56_io_out ? io_r_44_b : _GEN_22623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22625 = 9'h2d == r_count_56_io_out ? io_r_45_b : _GEN_22624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22626 = 9'h2e == r_count_56_io_out ? io_r_46_b : _GEN_22625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22627 = 9'h2f == r_count_56_io_out ? io_r_47_b : _GEN_22626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22628 = 9'h30 == r_count_56_io_out ? io_r_48_b : _GEN_22627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22629 = 9'h31 == r_count_56_io_out ? io_r_49_b : _GEN_22628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22630 = 9'h32 == r_count_56_io_out ? io_r_50_b : _GEN_22629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22631 = 9'h33 == r_count_56_io_out ? io_r_51_b : _GEN_22630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22632 = 9'h34 == r_count_56_io_out ? io_r_52_b : _GEN_22631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22633 = 9'h35 == r_count_56_io_out ? io_r_53_b : _GEN_22632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22634 = 9'h36 == r_count_56_io_out ? io_r_54_b : _GEN_22633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22635 = 9'h37 == r_count_56_io_out ? io_r_55_b : _GEN_22634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22636 = 9'h38 == r_count_56_io_out ? io_r_56_b : _GEN_22635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22637 = 9'h39 == r_count_56_io_out ? io_r_57_b : _GEN_22636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22638 = 9'h3a == r_count_56_io_out ? io_r_58_b : _GEN_22637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22639 = 9'h3b == r_count_56_io_out ? io_r_59_b : _GEN_22638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22640 = 9'h3c == r_count_56_io_out ? io_r_60_b : _GEN_22639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22641 = 9'h3d == r_count_56_io_out ? io_r_61_b : _GEN_22640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22642 = 9'h3e == r_count_56_io_out ? io_r_62_b : _GEN_22641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22643 = 9'h3f == r_count_56_io_out ? io_r_63_b : _GEN_22642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22644 = 9'h40 == r_count_56_io_out ? io_r_64_b : _GEN_22643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22645 = 9'h41 == r_count_56_io_out ? io_r_65_b : _GEN_22644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22646 = 9'h42 == r_count_56_io_out ? io_r_66_b : _GEN_22645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22647 = 9'h43 == r_count_56_io_out ? io_r_67_b : _GEN_22646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22648 = 9'h44 == r_count_56_io_out ? io_r_68_b : _GEN_22647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22649 = 9'h45 == r_count_56_io_out ? io_r_69_b : _GEN_22648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22650 = 9'h46 == r_count_56_io_out ? io_r_70_b : _GEN_22649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22651 = 9'h47 == r_count_56_io_out ? io_r_71_b : _GEN_22650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22652 = 9'h48 == r_count_56_io_out ? io_r_72_b : _GEN_22651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22653 = 9'h49 == r_count_56_io_out ? io_r_73_b : _GEN_22652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22654 = 9'h4a == r_count_56_io_out ? io_r_74_b : _GEN_22653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22655 = 9'h4b == r_count_56_io_out ? io_r_75_b : _GEN_22654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22656 = 9'h4c == r_count_56_io_out ? io_r_76_b : _GEN_22655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22657 = 9'h4d == r_count_56_io_out ? io_r_77_b : _GEN_22656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22658 = 9'h4e == r_count_56_io_out ? io_r_78_b : _GEN_22657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22659 = 9'h4f == r_count_56_io_out ? io_r_79_b : _GEN_22658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22660 = 9'h50 == r_count_56_io_out ? io_r_80_b : _GEN_22659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22661 = 9'h51 == r_count_56_io_out ? io_r_81_b : _GEN_22660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22662 = 9'h52 == r_count_56_io_out ? io_r_82_b : _GEN_22661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22663 = 9'h53 == r_count_56_io_out ? io_r_83_b : _GEN_22662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22664 = 9'h54 == r_count_56_io_out ? io_r_84_b : _GEN_22663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22665 = 9'h55 == r_count_56_io_out ? io_r_85_b : _GEN_22664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22666 = 9'h56 == r_count_56_io_out ? io_r_86_b : _GEN_22665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22667 = 9'h57 == r_count_56_io_out ? io_r_87_b : _GEN_22666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22668 = 9'h58 == r_count_56_io_out ? io_r_88_b : _GEN_22667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22669 = 9'h59 == r_count_56_io_out ? io_r_89_b : _GEN_22668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22670 = 9'h5a == r_count_56_io_out ? io_r_90_b : _GEN_22669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22671 = 9'h5b == r_count_56_io_out ? io_r_91_b : _GEN_22670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22672 = 9'h5c == r_count_56_io_out ? io_r_92_b : _GEN_22671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22673 = 9'h5d == r_count_56_io_out ? io_r_93_b : _GEN_22672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22674 = 9'h5e == r_count_56_io_out ? io_r_94_b : _GEN_22673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22675 = 9'h5f == r_count_56_io_out ? io_r_95_b : _GEN_22674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22676 = 9'h60 == r_count_56_io_out ? io_r_96_b : _GEN_22675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22677 = 9'h61 == r_count_56_io_out ? io_r_97_b : _GEN_22676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22678 = 9'h62 == r_count_56_io_out ? io_r_98_b : _GEN_22677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22679 = 9'h63 == r_count_56_io_out ? io_r_99_b : _GEN_22678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22680 = 9'h64 == r_count_56_io_out ? io_r_100_b : _GEN_22679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22681 = 9'h65 == r_count_56_io_out ? io_r_101_b : _GEN_22680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22682 = 9'h66 == r_count_56_io_out ? io_r_102_b : _GEN_22681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22683 = 9'h67 == r_count_56_io_out ? io_r_103_b : _GEN_22682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22684 = 9'h68 == r_count_56_io_out ? io_r_104_b : _GEN_22683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22685 = 9'h69 == r_count_56_io_out ? io_r_105_b : _GEN_22684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22686 = 9'h6a == r_count_56_io_out ? io_r_106_b : _GEN_22685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22687 = 9'h6b == r_count_56_io_out ? io_r_107_b : _GEN_22686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22688 = 9'h6c == r_count_56_io_out ? io_r_108_b : _GEN_22687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22689 = 9'h6d == r_count_56_io_out ? io_r_109_b : _GEN_22688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22690 = 9'h6e == r_count_56_io_out ? io_r_110_b : _GEN_22689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22691 = 9'h6f == r_count_56_io_out ? io_r_111_b : _GEN_22690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22692 = 9'h70 == r_count_56_io_out ? io_r_112_b : _GEN_22691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22693 = 9'h71 == r_count_56_io_out ? io_r_113_b : _GEN_22692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22694 = 9'h72 == r_count_56_io_out ? io_r_114_b : _GEN_22693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22695 = 9'h73 == r_count_56_io_out ? io_r_115_b : _GEN_22694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22696 = 9'h74 == r_count_56_io_out ? io_r_116_b : _GEN_22695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22697 = 9'h75 == r_count_56_io_out ? io_r_117_b : _GEN_22696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22698 = 9'h76 == r_count_56_io_out ? io_r_118_b : _GEN_22697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22699 = 9'h77 == r_count_56_io_out ? io_r_119_b : _GEN_22698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22700 = 9'h78 == r_count_56_io_out ? io_r_120_b : _GEN_22699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22701 = 9'h79 == r_count_56_io_out ? io_r_121_b : _GEN_22700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22702 = 9'h7a == r_count_56_io_out ? io_r_122_b : _GEN_22701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22703 = 9'h7b == r_count_56_io_out ? io_r_123_b : _GEN_22702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22704 = 9'h7c == r_count_56_io_out ? io_r_124_b : _GEN_22703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22705 = 9'h7d == r_count_56_io_out ? io_r_125_b : _GEN_22704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22706 = 9'h7e == r_count_56_io_out ? io_r_126_b : _GEN_22705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22707 = 9'h7f == r_count_56_io_out ? io_r_127_b : _GEN_22706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22708 = 9'h80 == r_count_56_io_out ? io_r_128_b : _GEN_22707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22709 = 9'h81 == r_count_56_io_out ? io_r_129_b : _GEN_22708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22710 = 9'h82 == r_count_56_io_out ? io_r_130_b : _GEN_22709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22711 = 9'h83 == r_count_56_io_out ? io_r_131_b : _GEN_22710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22712 = 9'h84 == r_count_56_io_out ? io_r_132_b : _GEN_22711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22713 = 9'h85 == r_count_56_io_out ? io_r_133_b : _GEN_22712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22714 = 9'h86 == r_count_56_io_out ? io_r_134_b : _GEN_22713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22715 = 9'h87 == r_count_56_io_out ? io_r_135_b : _GEN_22714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22716 = 9'h88 == r_count_56_io_out ? io_r_136_b : _GEN_22715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22717 = 9'h89 == r_count_56_io_out ? io_r_137_b : _GEN_22716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22718 = 9'h8a == r_count_56_io_out ? io_r_138_b : _GEN_22717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22719 = 9'h8b == r_count_56_io_out ? io_r_139_b : _GEN_22718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22720 = 9'h8c == r_count_56_io_out ? io_r_140_b : _GEN_22719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22721 = 9'h8d == r_count_56_io_out ? io_r_141_b : _GEN_22720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22722 = 9'h8e == r_count_56_io_out ? io_r_142_b : _GEN_22721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22723 = 9'h8f == r_count_56_io_out ? io_r_143_b : _GEN_22722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22724 = 9'h90 == r_count_56_io_out ? io_r_144_b : _GEN_22723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22725 = 9'h91 == r_count_56_io_out ? io_r_145_b : _GEN_22724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22726 = 9'h92 == r_count_56_io_out ? io_r_146_b : _GEN_22725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22727 = 9'h93 == r_count_56_io_out ? io_r_147_b : _GEN_22726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22728 = 9'h94 == r_count_56_io_out ? io_r_148_b : _GEN_22727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22729 = 9'h95 == r_count_56_io_out ? io_r_149_b : _GEN_22728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22730 = 9'h96 == r_count_56_io_out ? io_r_150_b : _GEN_22729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22731 = 9'h97 == r_count_56_io_out ? io_r_151_b : _GEN_22730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22732 = 9'h98 == r_count_56_io_out ? io_r_152_b : _GEN_22731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22733 = 9'h99 == r_count_56_io_out ? io_r_153_b : _GEN_22732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22734 = 9'h9a == r_count_56_io_out ? io_r_154_b : _GEN_22733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22735 = 9'h9b == r_count_56_io_out ? io_r_155_b : _GEN_22734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22736 = 9'h9c == r_count_56_io_out ? io_r_156_b : _GEN_22735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22737 = 9'h9d == r_count_56_io_out ? io_r_157_b : _GEN_22736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22738 = 9'h9e == r_count_56_io_out ? io_r_158_b : _GEN_22737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22739 = 9'h9f == r_count_56_io_out ? io_r_159_b : _GEN_22738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22740 = 9'ha0 == r_count_56_io_out ? io_r_160_b : _GEN_22739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22741 = 9'ha1 == r_count_56_io_out ? io_r_161_b : _GEN_22740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22742 = 9'ha2 == r_count_56_io_out ? io_r_162_b : _GEN_22741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22743 = 9'ha3 == r_count_56_io_out ? io_r_163_b : _GEN_22742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22744 = 9'ha4 == r_count_56_io_out ? io_r_164_b : _GEN_22743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22745 = 9'ha5 == r_count_56_io_out ? io_r_165_b : _GEN_22744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22746 = 9'ha6 == r_count_56_io_out ? io_r_166_b : _GEN_22745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22747 = 9'ha7 == r_count_56_io_out ? io_r_167_b : _GEN_22746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22748 = 9'ha8 == r_count_56_io_out ? io_r_168_b : _GEN_22747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22749 = 9'ha9 == r_count_56_io_out ? io_r_169_b : _GEN_22748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22750 = 9'haa == r_count_56_io_out ? io_r_170_b : _GEN_22749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22751 = 9'hab == r_count_56_io_out ? io_r_171_b : _GEN_22750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22752 = 9'hac == r_count_56_io_out ? io_r_172_b : _GEN_22751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22753 = 9'had == r_count_56_io_out ? io_r_173_b : _GEN_22752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22754 = 9'hae == r_count_56_io_out ? io_r_174_b : _GEN_22753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22755 = 9'haf == r_count_56_io_out ? io_r_175_b : _GEN_22754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22756 = 9'hb0 == r_count_56_io_out ? io_r_176_b : _GEN_22755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22757 = 9'hb1 == r_count_56_io_out ? io_r_177_b : _GEN_22756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22758 = 9'hb2 == r_count_56_io_out ? io_r_178_b : _GEN_22757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22759 = 9'hb3 == r_count_56_io_out ? io_r_179_b : _GEN_22758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22760 = 9'hb4 == r_count_56_io_out ? io_r_180_b : _GEN_22759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22761 = 9'hb5 == r_count_56_io_out ? io_r_181_b : _GEN_22760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22762 = 9'hb6 == r_count_56_io_out ? io_r_182_b : _GEN_22761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22763 = 9'hb7 == r_count_56_io_out ? io_r_183_b : _GEN_22762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22764 = 9'hb8 == r_count_56_io_out ? io_r_184_b : _GEN_22763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22765 = 9'hb9 == r_count_56_io_out ? io_r_185_b : _GEN_22764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22766 = 9'hba == r_count_56_io_out ? io_r_186_b : _GEN_22765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22767 = 9'hbb == r_count_56_io_out ? io_r_187_b : _GEN_22766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22768 = 9'hbc == r_count_56_io_out ? io_r_188_b : _GEN_22767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22769 = 9'hbd == r_count_56_io_out ? io_r_189_b : _GEN_22768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22770 = 9'hbe == r_count_56_io_out ? io_r_190_b : _GEN_22769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22771 = 9'hbf == r_count_56_io_out ? io_r_191_b : _GEN_22770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22772 = 9'hc0 == r_count_56_io_out ? io_r_192_b : _GEN_22771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22773 = 9'hc1 == r_count_56_io_out ? io_r_193_b : _GEN_22772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22774 = 9'hc2 == r_count_56_io_out ? io_r_194_b : _GEN_22773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22775 = 9'hc3 == r_count_56_io_out ? io_r_195_b : _GEN_22774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22776 = 9'hc4 == r_count_56_io_out ? io_r_196_b : _GEN_22775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22777 = 9'hc5 == r_count_56_io_out ? io_r_197_b : _GEN_22776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22778 = 9'hc6 == r_count_56_io_out ? io_r_198_b : _GEN_22777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22779 = 9'hc7 == r_count_56_io_out ? io_r_199_b : _GEN_22778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22780 = 9'hc8 == r_count_56_io_out ? io_r_200_b : _GEN_22779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22781 = 9'hc9 == r_count_56_io_out ? io_r_201_b : _GEN_22780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22782 = 9'hca == r_count_56_io_out ? io_r_202_b : _GEN_22781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22783 = 9'hcb == r_count_56_io_out ? io_r_203_b : _GEN_22782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22784 = 9'hcc == r_count_56_io_out ? io_r_204_b : _GEN_22783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22785 = 9'hcd == r_count_56_io_out ? io_r_205_b : _GEN_22784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22786 = 9'hce == r_count_56_io_out ? io_r_206_b : _GEN_22785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22787 = 9'hcf == r_count_56_io_out ? io_r_207_b : _GEN_22786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22788 = 9'hd0 == r_count_56_io_out ? io_r_208_b : _GEN_22787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22789 = 9'hd1 == r_count_56_io_out ? io_r_209_b : _GEN_22788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22790 = 9'hd2 == r_count_56_io_out ? io_r_210_b : _GEN_22789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22791 = 9'hd3 == r_count_56_io_out ? io_r_211_b : _GEN_22790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22792 = 9'hd4 == r_count_56_io_out ? io_r_212_b : _GEN_22791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22793 = 9'hd5 == r_count_56_io_out ? io_r_213_b : _GEN_22792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22794 = 9'hd6 == r_count_56_io_out ? io_r_214_b : _GEN_22793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22795 = 9'hd7 == r_count_56_io_out ? io_r_215_b : _GEN_22794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22796 = 9'hd8 == r_count_56_io_out ? io_r_216_b : _GEN_22795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22797 = 9'hd9 == r_count_56_io_out ? io_r_217_b : _GEN_22796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22798 = 9'hda == r_count_56_io_out ? io_r_218_b : _GEN_22797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22799 = 9'hdb == r_count_56_io_out ? io_r_219_b : _GEN_22798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22800 = 9'hdc == r_count_56_io_out ? io_r_220_b : _GEN_22799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22801 = 9'hdd == r_count_56_io_out ? io_r_221_b : _GEN_22800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22802 = 9'hde == r_count_56_io_out ? io_r_222_b : _GEN_22801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22803 = 9'hdf == r_count_56_io_out ? io_r_223_b : _GEN_22802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22804 = 9'he0 == r_count_56_io_out ? io_r_224_b : _GEN_22803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22805 = 9'he1 == r_count_56_io_out ? io_r_225_b : _GEN_22804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22806 = 9'he2 == r_count_56_io_out ? io_r_226_b : _GEN_22805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22807 = 9'he3 == r_count_56_io_out ? io_r_227_b : _GEN_22806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22808 = 9'he4 == r_count_56_io_out ? io_r_228_b : _GEN_22807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22809 = 9'he5 == r_count_56_io_out ? io_r_229_b : _GEN_22808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22810 = 9'he6 == r_count_56_io_out ? io_r_230_b : _GEN_22809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22811 = 9'he7 == r_count_56_io_out ? io_r_231_b : _GEN_22810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22812 = 9'he8 == r_count_56_io_out ? io_r_232_b : _GEN_22811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22813 = 9'he9 == r_count_56_io_out ? io_r_233_b : _GEN_22812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22814 = 9'hea == r_count_56_io_out ? io_r_234_b : _GEN_22813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22815 = 9'heb == r_count_56_io_out ? io_r_235_b : _GEN_22814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22816 = 9'hec == r_count_56_io_out ? io_r_236_b : _GEN_22815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22817 = 9'hed == r_count_56_io_out ? io_r_237_b : _GEN_22816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22818 = 9'hee == r_count_56_io_out ? io_r_238_b : _GEN_22817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22819 = 9'hef == r_count_56_io_out ? io_r_239_b : _GEN_22818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22820 = 9'hf0 == r_count_56_io_out ? io_r_240_b : _GEN_22819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22821 = 9'hf1 == r_count_56_io_out ? io_r_241_b : _GEN_22820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22822 = 9'hf2 == r_count_56_io_out ? io_r_242_b : _GEN_22821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22823 = 9'hf3 == r_count_56_io_out ? io_r_243_b : _GEN_22822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22824 = 9'hf4 == r_count_56_io_out ? io_r_244_b : _GEN_22823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22825 = 9'hf5 == r_count_56_io_out ? io_r_245_b : _GEN_22824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22826 = 9'hf6 == r_count_56_io_out ? io_r_246_b : _GEN_22825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22827 = 9'hf7 == r_count_56_io_out ? io_r_247_b : _GEN_22826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22828 = 9'hf8 == r_count_56_io_out ? io_r_248_b : _GEN_22827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22829 = 9'hf9 == r_count_56_io_out ? io_r_249_b : _GEN_22828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22830 = 9'hfa == r_count_56_io_out ? io_r_250_b : _GEN_22829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22831 = 9'hfb == r_count_56_io_out ? io_r_251_b : _GEN_22830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22832 = 9'hfc == r_count_56_io_out ? io_r_252_b : _GEN_22831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22833 = 9'hfd == r_count_56_io_out ? io_r_253_b : _GEN_22832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22834 = 9'hfe == r_count_56_io_out ? io_r_254_b : _GEN_22833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22835 = 9'hff == r_count_56_io_out ? io_r_255_b : _GEN_22834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22836 = 9'h100 == r_count_56_io_out ? io_r_256_b : _GEN_22835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22837 = 9'h101 == r_count_56_io_out ? io_r_257_b : _GEN_22836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22838 = 9'h102 == r_count_56_io_out ? io_r_258_b : _GEN_22837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22839 = 9'h103 == r_count_56_io_out ? io_r_259_b : _GEN_22838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22840 = 9'h104 == r_count_56_io_out ? io_r_260_b : _GEN_22839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22841 = 9'h105 == r_count_56_io_out ? io_r_261_b : _GEN_22840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22842 = 9'h106 == r_count_56_io_out ? io_r_262_b : _GEN_22841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22843 = 9'h107 == r_count_56_io_out ? io_r_263_b : _GEN_22842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22844 = 9'h108 == r_count_56_io_out ? io_r_264_b : _GEN_22843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22845 = 9'h109 == r_count_56_io_out ? io_r_265_b : _GEN_22844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22846 = 9'h10a == r_count_56_io_out ? io_r_266_b : _GEN_22845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22847 = 9'h10b == r_count_56_io_out ? io_r_267_b : _GEN_22846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22848 = 9'h10c == r_count_56_io_out ? io_r_268_b : _GEN_22847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22849 = 9'h10d == r_count_56_io_out ? io_r_269_b : _GEN_22848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22850 = 9'h10e == r_count_56_io_out ? io_r_270_b : _GEN_22849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22851 = 9'h10f == r_count_56_io_out ? io_r_271_b : _GEN_22850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22852 = 9'h110 == r_count_56_io_out ? io_r_272_b : _GEN_22851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22853 = 9'h111 == r_count_56_io_out ? io_r_273_b : _GEN_22852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22854 = 9'h112 == r_count_56_io_out ? io_r_274_b : _GEN_22853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22855 = 9'h113 == r_count_56_io_out ? io_r_275_b : _GEN_22854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22856 = 9'h114 == r_count_56_io_out ? io_r_276_b : _GEN_22855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22857 = 9'h115 == r_count_56_io_out ? io_r_277_b : _GEN_22856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22858 = 9'h116 == r_count_56_io_out ? io_r_278_b : _GEN_22857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22859 = 9'h117 == r_count_56_io_out ? io_r_279_b : _GEN_22858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22860 = 9'h118 == r_count_56_io_out ? io_r_280_b : _GEN_22859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22861 = 9'h119 == r_count_56_io_out ? io_r_281_b : _GEN_22860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22862 = 9'h11a == r_count_56_io_out ? io_r_282_b : _GEN_22861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22863 = 9'h11b == r_count_56_io_out ? io_r_283_b : _GEN_22862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22864 = 9'h11c == r_count_56_io_out ? io_r_284_b : _GEN_22863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22865 = 9'h11d == r_count_56_io_out ? io_r_285_b : _GEN_22864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22866 = 9'h11e == r_count_56_io_out ? io_r_286_b : _GEN_22865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22867 = 9'h11f == r_count_56_io_out ? io_r_287_b : _GEN_22866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22868 = 9'h120 == r_count_56_io_out ? io_r_288_b : _GEN_22867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22869 = 9'h121 == r_count_56_io_out ? io_r_289_b : _GEN_22868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22870 = 9'h122 == r_count_56_io_out ? io_r_290_b : _GEN_22869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22871 = 9'h123 == r_count_56_io_out ? io_r_291_b : _GEN_22870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22872 = 9'h124 == r_count_56_io_out ? io_r_292_b : _GEN_22871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22873 = 9'h125 == r_count_56_io_out ? io_r_293_b : _GEN_22872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22874 = 9'h126 == r_count_56_io_out ? io_r_294_b : _GEN_22873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22875 = 9'h127 == r_count_56_io_out ? io_r_295_b : _GEN_22874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22876 = 9'h128 == r_count_56_io_out ? io_r_296_b : _GEN_22875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22877 = 9'h129 == r_count_56_io_out ? io_r_297_b : _GEN_22876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22878 = 9'h12a == r_count_56_io_out ? io_r_298_b : _GEN_22877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22879 = 9'h12b == r_count_56_io_out ? io_r_299_b : _GEN_22878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22880 = 9'h12c == r_count_56_io_out ? io_r_300_b : _GEN_22879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22881 = 9'h12d == r_count_56_io_out ? io_r_301_b : _GEN_22880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22882 = 9'h12e == r_count_56_io_out ? io_r_302_b : _GEN_22881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22883 = 9'h12f == r_count_56_io_out ? io_r_303_b : _GEN_22882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22884 = 9'h130 == r_count_56_io_out ? io_r_304_b : _GEN_22883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22885 = 9'h131 == r_count_56_io_out ? io_r_305_b : _GEN_22884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22886 = 9'h132 == r_count_56_io_out ? io_r_306_b : _GEN_22885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22887 = 9'h133 == r_count_56_io_out ? io_r_307_b : _GEN_22886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22888 = 9'h134 == r_count_56_io_out ? io_r_308_b : _GEN_22887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22889 = 9'h135 == r_count_56_io_out ? io_r_309_b : _GEN_22888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22890 = 9'h136 == r_count_56_io_out ? io_r_310_b : _GEN_22889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22891 = 9'h137 == r_count_56_io_out ? io_r_311_b : _GEN_22890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22892 = 9'h138 == r_count_56_io_out ? io_r_312_b : _GEN_22891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22893 = 9'h139 == r_count_56_io_out ? io_r_313_b : _GEN_22892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22894 = 9'h13a == r_count_56_io_out ? io_r_314_b : _GEN_22893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22895 = 9'h13b == r_count_56_io_out ? io_r_315_b : _GEN_22894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22896 = 9'h13c == r_count_56_io_out ? io_r_316_b : _GEN_22895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22897 = 9'h13d == r_count_56_io_out ? io_r_317_b : _GEN_22896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22898 = 9'h13e == r_count_56_io_out ? io_r_318_b : _GEN_22897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22899 = 9'h13f == r_count_56_io_out ? io_r_319_b : _GEN_22898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22900 = 9'h140 == r_count_56_io_out ? io_r_320_b : _GEN_22899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22901 = 9'h141 == r_count_56_io_out ? io_r_321_b : _GEN_22900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22902 = 9'h142 == r_count_56_io_out ? io_r_322_b : _GEN_22901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22903 = 9'h143 == r_count_56_io_out ? io_r_323_b : _GEN_22902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22904 = 9'h144 == r_count_56_io_out ? io_r_324_b : _GEN_22903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22905 = 9'h145 == r_count_56_io_out ? io_r_325_b : _GEN_22904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22906 = 9'h146 == r_count_56_io_out ? io_r_326_b : _GEN_22905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22907 = 9'h147 == r_count_56_io_out ? io_r_327_b : _GEN_22906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22908 = 9'h148 == r_count_56_io_out ? io_r_328_b : _GEN_22907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22909 = 9'h149 == r_count_56_io_out ? io_r_329_b : _GEN_22908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22910 = 9'h14a == r_count_56_io_out ? io_r_330_b : _GEN_22909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22911 = 9'h14b == r_count_56_io_out ? io_r_331_b : _GEN_22910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22912 = 9'h14c == r_count_56_io_out ? io_r_332_b : _GEN_22911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22913 = 9'h14d == r_count_56_io_out ? io_r_333_b : _GEN_22912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22914 = 9'h14e == r_count_56_io_out ? io_r_334_b : _GEN_22913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22915 = 9'h14f == r_count_56_io_out ? io_r_335_b : _GEN_22914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22916 = 9'h150 == r_count_56_io_out ? io_r_336_b : _GEN_22915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22917 = 9'h151 == r_count_56_io_out ? io_r_337_b : _GEN_22916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22918 = 9'h152 == r_count_56_io_out ? io_r_338_b : _GEN_22917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22919 = 9'h153 == r_count_56_io_out ? io_r_339_b : _GEN_22918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22920 = 9'h154 == r_count_56_io_out ? io_r_340_b : _GEN_22919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22921 = 9'h155 == r_count_56_io_out ? io_r_341_b : _GEN_22920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22922 = 9'h156 == r_count_56_io_out ? io_r_342_b : _GEN_22921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22923 = 9'h157 == r_count_56_io_out ? io_r_343_b : _GEN_22922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22924 = 9'h158 == r_count_56_io_out ? io_r_344_b : _GEN_22923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22925 = 9'h159 == r_count_56_io_out ? io_r_345_b : _GEN_22924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22926 = 9'h15a == r_count_56_io_out ? io_r_346_b : _GEN_22925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22927 = 9'h15b == r_count_56_io_out ? io_r_347_b : _GEN_22926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22928 = 9'h15c == r_count_56_io_out ? io_r_348_b : _GEN_22927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22929 = 9'h15d == r_count_56_io_out ? io_r_349_b : _GEN_22928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22930 = 9'h15e == r_count_56_io_out ? io_r_350_b : _GEN_22929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22931 = 9'h15f == r_count_56_io_out ? io_r_351_b : _GEN_22930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22932 = 9'h160 == r_count_56_io_out ? io_r_352_b : _GEN_22931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22933 = 9'h161 == r_count_56_io_out ? io_r_353_b : _GEN_22932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22934 = 9'h162 == r_count_56_io_out ? io_r_354_b : _GEN_22933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22935 = 9'h163 == r_count_56_io_out ? io_r_355_b : _GEN_22934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22936 = 9'h164 == r_count_56_io_out ? io_r_356_b : _GEN_22935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22937 = 9'h165 == r_count_56_io_out ? io_r_357_b : _GEN_22936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22938 = 9'h166 == r_count_56_io_out ? io_r_358_b : _GEN_22937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22939 = 9'h167 == r_count_56_io_out ? io_r_359_b : _GEN_22938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22940 = 9'h168 == r_count_56_io_out ? io_r_360_b : _GEN_22939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22941 = 9'h169 == r_count_56_io_out ? io_r_361_b : _GEN_22940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22942 = 9'h16a == r_count_56_io_out ? io_r_362_b : _GEN_22941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22943 = 9'h16b == r_count_56_io_out ? io_r_363_b : _GEN_22942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22944 = 9'h16c == r_count_56_io_out ? io_r_364_b : _GEN_22943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22945 = 9'h16d == r_count_56_io_out ? io_r_365_b : _GEN_22944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22946 = 9'h16e == r_count_56_io_out ? io_r_366_b : _GEN_22945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22947 = 9'h16f == r_count_56_io_out ? io_r_367_b : _GEN_22946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22948 = 9'h170 == r_count_56_io_out ? io_r_368_b : _GEN_22947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22949 = 9'h171 == r_count_56_io_out ? io_r_369_b : _GEN_22948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22950 = 9'h172 == r_count_56_io_out ? io_r_370_b : _GEN_22949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22951 = 9'h173 == r_count_56_io_out ? io_r_371_b : _GEN_22950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22952 = 9'h174 == r_count_56_io_out ? io_r_372_b : _GEN_22951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22953 = 9'h175 == r_count_56_io_out ? io_r_373_b : _GEN_22952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22954 = 9'h176 == r_count_56_io_out ? io_r_374_b : _GEN_22953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22955 = 9'h177 == r_count_56_io_out ? io_r_375_b : _GEN_22954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22956 = 9'h178 == r_count_56_io_out ? io_r_376_b : _GEN_22955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22957 = 9'h179 == r_count_56_io_out ? io_r_377_b : _GEN_22956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22958 = 9'h17a == r_count_56_io_out ? io_r_378_b : _GEN_22957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22959 = 9'h17b == r_count_56_io_out ? io_r_379_b : _GEN_22958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22960 = 9'h17c == r_count_56_io_out ? io_r_380_b : _GEN_22959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22961 = 9'h17d == r_count_56_io_out ? io_r_381_b : _GEN_22960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22962 = 9'h17e == r_count_56_io_out ? io_r_382_b : _GEN_22961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22963 = 9'h17f == r_count_56_io_out ? io_r_383_b : _GEN_22962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22964 = 9'h180 == r_count_56_io_out ? io_r_384_b : _GEN_22963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22965 = 9'h181 == r_count_56_io_out ? io_r_385_b : _GEN_22964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22966 = 9'h182 == r_count_56_io_out ? io_r_386_b : _GEN_22965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22967 = 9'h183 == r_count_56_io_out ? io_r_387_b : _GEN_22966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22968 = 9'h184 == r_count_56_io_out ? io_r_388_b : _GEN_22967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22969 = 9'h185 == r_count_56_io_out ? io_r_389_b : _GEN_22968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22970 = 9'h186 == r_count_56_io_out ? io_r_390_b : _GEN_22969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22971 = 9'h187 == r_count_56_io_out ? io_r_391_b : _GEN_22970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22972 = 9'h188 == r_count_56_io_out ? io_r_392_b : _GEN_22971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22973 = 9'h189 == r_count_56_io_out ? io_r_393_b : _GEN_22972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22974 = 9'h18a == r_count_56_io_out ? io_r_394_b : _GEN_22973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22975 = 9'h18b == r_count_56_io_out ? io_r_395_b : _GEN_22974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22976 = 9'h18c == r_count_56_io_out ? io_r_396_b : _GEN_22975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22977 = 9'h18d == r_count_56_io_out ? io_r_397_b : _GEN_22976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22978 = 9'h18e == r_count_56_io_out ? io_r_398_b : _GEN_22977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22981 = 9'h1 == r_count_57_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22982 = 9'h2 == r_count_57_io_out ? io_r_2_b : _GEN_22981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22983 = 9'h3 == r_count_57_io_out ? io_r_3_b : _GEN_22982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22984 = 9'h4 == r_count_57_io_out ? io_r_4_b : _GEN_22983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22985 = 9'h5 == r_count_57_io_out ? io_r_5_b : _GEN_22984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22986 = 9'h6 == r_count_57_io_out ? io_r_6_b : _GEN_22985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22987 = 9'h7 == r_count_57_io_out ? io_r_7_b : _GEN_22986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22988 = 9'h8 == r_count_57_io_out ? io_r_8_b : _GEN_22987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22989 = 9'h9 == r_count_57_io_out ? io_r_9_b : _GEN_22988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22990 = 9'ha == r_count_57_io_out ? io_r_10_b : _GEN_22989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22991 = 9'hb == r_count_57_io_out ? io_r_11_b : _GEN_22990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22992 = 9'hc == r_count_57_io_out ? io_r_12_b : _GEN_22991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22993 = 9'hd == r_count_57_io_out ? io_r_13_b : _GEN_22992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22994 = 9'he == r_count_57_io_out ? io_r_14_b : _GEN_22993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22995 = 9'hf == r_count_57_io_out ? io_r_15_b : _GEN_22994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22996 = 9'h10 == r_count_57_io_out ? io_r_16_b : _GEN_22995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22997 = 9'h11 == r_count_57_io_out ? io_r_17_b : _GEN_22996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22998 = 9'h12 == r_count_57_io_out ? io_r_18_b : _GEN_22997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22999 = 9'h13 == r_count_57_io_out ? io_r_19_b : _GEN_22998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23000 = 9'h14 == r_count_57_io_out ? io_r_20_b : _GEN_22999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23001 = 9'h15 == r_count_57_io_out ? io_r_21_b : _GEN_23000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23002 = 9'h16 == r_count_57_io_out ? io_r_22_b : _GEN_23001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23003 = 9'h17 == r_count_57_io_out ? io_r_23_b : _GEN_23002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23004 = 9'h18 == r_count_57_io_out ? io_r_24_b : _GEN_23003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23005 = 9'h19 == r_count_57_io_out ? io_r_25_b : _GEN_23004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23006 = 9'h1a == r_count_57_io_out ? io_r_26_b : _GEN_23005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23007 = 9'h1b == r_count_57_io_out ? io_r_27_b : _GEN_23006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23008 = 9'h1c == r_count_57_io_out ? io_r_28_b : _GEN_23007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23009 = 9'h1d == r_count_57_io_out ? io_r_29_b : _GEN_23008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23010 = 9'h1e == r_count_57_io_out ? io_r_30_b : _GEN_23009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23011 = 9'h1f == r_count_57_io_out ? io_r_31_b : _GEN_23010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23012 = 9'h20 == r_count_57_io_out ? io_r_32_b : _GEN_23011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23013 = 9'h21 == r_count_57_io_out ? io_r_33_b : _GEN_23012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23014 = 9'h22 == r_count_57_io_out ? io_r_34_b : _GEN_23013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23015 = 9'h23 == r_count_57_io_out ? io_r_35_b : _GEN_23014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23016 = 9'h24 == r_count_57_io_out ? io_r_36_b : _GEN_23015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23017 = 9'h25 == r_count_57_io_out ? io_r_37_b : _GEN_23016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23018 = 9'h26 == r_count_57_io_out ? io_r_38_b : _GEN_23017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23019 = 9'h27 == r_count_57_io_out ? io_r_39_b : _GEN_23018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23020 = 9'h28 == r_count_57_io_out ? io_r_40_b : _GEN_23019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23021 = 9'h29 == r_count_57_io_out ? io_r_41_b : _GEN_23020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23022 = 9'h2a == r_count_57_io_out ? io_r_42_b : _GEN_23021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23023 = 9'h2b == r_count_57_io_out ? io_r_43_b : _GEN_23022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23024 = 9'h2c == r_count_57_io_out ? io_r_44_b : _GEN_23023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23025 = 9'h2d == r_count_57_io_out ? io_r_45_b : _GEN_23024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23026 = 9'h2e == r_count_57_io_out ? io_r_46_b : _GEN_23025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23027 = 9'h2f == r_count_57_io_out ? io_r_47_b : _GEN_23026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23028 = 9'h30 == r_count_57_io_out ? io_r_48_b : _GEN_23027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23029 = 9'h31 == r_count_57_io_out ? io_r_49_b : _GEN_23028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23030 = 9'h32 == r_count_57_io_out ? io_r_50_b : _GEN_23029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23031 = 9'h33 == r_count_57_io_out ? io_r_51_b : _GEN_23030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23032 = 9'h34 == r_count_57_io_out ? io_r_52_b : _GEN_23031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23033 = 9'h35 == r_count_57_io_out ? io_r_53_b : _GEN_23032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23034 = 9'h36 == r_count_57_io_out ? io_r_54_b : _GEN_23033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23035 = 9'h37 == r_count_57_io_out ? io_r_55_b : _GEN_23034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23036 = 9'h38 == r_count_57_io_out ? io_r_56_b : _GEN_23035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23037 = 9'h39 == r_count_57_io_out ? io_r_57_b : _GEN_23036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23038 = 9'h3a == r_count_57_io_out ? io_r_58_b : _GEN_23037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23039 = 9'h3b == r_count_57_io_out ? io_r_59_b : _GEN_23038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23040 = 9'h3c == r_count_57_io_out ? io_r_60_b : _GEN_23039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23041 = 9'h3d == r_count_57_io_out ? io_r_61_b : _GEN_23040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23042 = 9'h3e == r_count_57_io_out ? io_r_62_b : _GEN_23041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23043 = 9'h3f == r_count_57_io_out ? io_r_63_b : _GEN_23042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23044 = 9'h40 == r_count_57_io_out ? io_r_64_b : _GEN_23043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23045 = 9'h41 == r_count_57_io_out ? io_r_65_b : _GEN_23044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23046 = 9'h42 == r_count_57_io_out ? io_r_66_b : _GEN_23045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23047 = 9'h43 == r_count_57_io_out ? io_r_67_b : _GEN_23046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23048 = 9'h44 == r_count_57_io_out ? io_r_68_b : _GEN_23047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23049 = 9'h45 == r_count_57_io_out ? io_r_69_b : _GEN_23048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23050 = 9'h46 == r_count_57_io_out ? io_r_70_b : _GEN_23049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23051 = 9'h47 == r_count_57_io_out ? io_r_71_b : _GEN_23050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23052 = 9'h48 == r_count_57_io_out ? io_r_72_b : _GEN_23051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23053 = 9'h49 == r_count_57_io_out ? io_r_73_b : _GEN_23052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23054 = 9'h4a == r_count_57_io_out ? io_r_74_b : _GEN_23053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23055 = 9'h4b == r_count_57_io_out ? io_r_75_b : _GEN_23054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23056 = 9'h4c == r_count_57_io_out ? io_r_76_b : _GEN_23055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23057 = 9'h4d == r_count_57_io_out ? io_r_77_b : _GEN_23056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23058 = 9'h4e == r_count_57_io_out ? io_r_78_b : _GEN_23057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23059 = 9'h4f == r_count_57_io_out ? io_r_79_b : _GEN_23058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23060 = 9'h50 == r_count_57_io_out ? io_r_80_b : _GEN_23059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23061 = 9'h51 == r_count_57_io_out ? io_r_81_b : _GEN_23060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23062 = 9'h52 == r_count_57_io_out ? io_r_82_b : _GEN_23061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23063 = 9'h53 == r_count_57_io_out ? io_r_83_b : _GEN_23062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23064 = 9'h54 == r_count_57_io_out ? io_r_84_b : _GEN_23063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23065 = 9'h55 == r_count_57_io_out ? io_r_85_b : _GEN_23064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23066 = 9'h56 == r_count_57_io_out ? io_r_86_b : _GEN_23065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23067 = 9'h57 == r_count_57_io_out ? io_r_87_b : _GEN_23066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23068 = 9'h58 == r_count_57_io_out ? io_r_88_b : _GEN_23067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23069 = 9'h59 == r_count_57_io_out ? io_r_89_b : _GEN_23068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23070 = 9'h5a == r_count_57_io_out ? io_r_90_b : _GEN_23069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23071 = 9'h5b == r_count_57_io_out ? io_r_91_b : _GEN_23070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23072 = 9'h5c == r_count_57_io_out ? io_r_92_b : _GEN_23071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23073 = 9'h5d == r_count_57_io_out ? io_r_93_b : _GEN_23072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23074 = 9'h5e == r_count_57_io_out ? io_r_94_b : _GEN_23073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23075 = 9'h5f == r_count_57_io_out ? io_r_95_b : _GEN_23074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23076 = 9'h60 == r_count_57_io_out ? io_r_96_b : _GEN_23075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23077 = 9'h61 == r_count_57_io_out ? io_r_97_b : _GEN_23076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23078 = 9'h62 == r_count_57_io_out ? io_r_98_b : _GEN_23077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23079 = 9'h63 == r_count_57_io_out ? io_r_99_b : _GEN_23078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23080 = 9'h64 == r_count_57_io_out ? io_r_100_b : _GEN_23079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23081 = 9'h65 == r_count_57_io_out ? io_r_101_b : _GEN_23080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23082 = 9'h66 == r_count_57_io_out ? io_r_102_b : _GEN_23081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23083 = 9'h67 == r_count_57_io_out ? io_r_103_b : _GEN_23082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23084 = 9'h68 == r_count_57_io_out ? io_r_104_b : _GEN_23083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23085 = 9'h69 == r_count_57_io_out ? io_r_105_b : _GEN_23084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23086 = 9'h6a == r_count_57_io_out ? io_r_106_b : _GEN_23085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23087 = 9'h6b == r_count_57_io_out ? io_r_107_b : _GEN_23086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23088 = 9'h6c == r_count_57_io_out ? io_r_108_b : _GEN_23087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23089 = 9'h6d == r_count_57_io_out ? io_r_109_b : _GEN_23088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23090 = 9'h6e == r_count_57_io_out ? io_r_110_b : _GEN_23089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23091 = 9'h6f == r_count_57_io_out ? io_r_111_b : _GEN_23090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23092 = 9'h70 == r_count_57_io_out ? io_r_112_b : _GEN_23091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23093 = 9'h71 == r_count_57_io_out ? io_r_113_b : _GEN_23092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23094 = 9'h72 == r_count_57_io_out ? io_r_114_b : _GEN_23093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23095 = 9'h73 == r_count_57_io_out ? io_r_115_b : _GEN_23094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23096 = 9'h74 == r_count_57_io_out ? io_r_116_b : _GEN_23095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23097 = 9'h75 == r_count_57_io_out ? io_r_117_b : _GEN_23096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23098 = 9'h76 == r_count_57_io_out ? io_r_118_b : _GEN_23097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23099 = 9'h77 == r_count_57_io_out ? io_r_119_b : _GEN_23098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23100 = 9'h78 == r_count_57_io_out ? io_r_120_b : _GEN_23099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23101 = 9'h79 == r_count_57_io_out ? io_r_121_b : _GEN_23100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23102 = 9'h7a == r_count_57_io_out ? io_r_122_b : _GEN_23101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23103 = 9'h7b == r_count_57_io_out ? io_r_123_b : _GEN_23102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23104 = 9'h7c == r_count_57_io_out ? io_r_124_b : _GEN_23103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23105 = 9'h7d == r_count_57_io_out ? io_r_125_b : _GEN_23104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23106 = 9'h7e == r_count_57_io_out ? io_r_126_b : _GEN_23105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23107 = 9'h7f == r_count_57_io_out ? io_r_127_b : _GEN_23106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23108 = 9'h80 == r_count_57_io_out ? io_r_128_b : _GEN_23107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23109 = 9'h81 == r_count_57_io_out ? io_r_129_b : _GEN_23108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23110 = 9'h82 == r_count_57_io_out ? io_r_130_b : _GEN_23109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23111 = 9'h83 == r_count_57_io_out ? io_r_131_b : _GEN_23110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23112 = 9'h84 == r_count_57_io_out ? io_r_132_b : _GEN_23111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23113 = 9'h85 == r_count_57_io_out ? io_r_133_b : _GEN_23112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23114 = 9'h86 == r_count_57_io_out ? io_r_134_b : _GEN_23113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23115 = 9'h87 == r_count_57_io_out ? io_r_135_b : _GEN_23114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23116 = 9'h88 == r_count_57_io_out ? io_r_136_b : _GEN_23115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23117 = 9'h89 == r_count_57_io_out ? io_r_137_b : _GEN_23116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23118 = 9'h8a == r_count_57_io_out ? io_r_138_b : _GEN_23117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23119 = 9'h8b == r_count_57_io_out ? io_r_139_b : _GEN_23118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23120 = 9'h8c == r_count_57_io_out ? io_r_140_b : _GEN_23119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23121 = 9'h8d == r_count_57_io_out ? io_r_141_b : _GEN_23120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23122 = 9'h8e == r_count_57_io_out ? io_r_142_b : _GEN_23121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23123 = 9'h8f == r_count_57_io_out ? io_r_143_b : _GEN_23122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23124 = 9'h90 == r_count_57_io_out ? io_r_144_b : _GEN_23123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23125 = 9'h91 == r_count_57_io_out ? io_r_145_b : _GEN_23124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23126 = 9'h92 == r_count_57_io_out ? io_r_146_b : _GEN_23125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23127 = 9'h93 == r_count_57_io_out ? io_r_147_b : _GEN_23126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23128 = 9'h94 == r_count_57_io_out ? io_r_148_b : _GEN_23127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23129 = 9'h95 == r_count_57_io_out ? io_r_149_b : _GEN_23128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23130 = 9'h96 == r_count_57_io_out ? io_r_150_b : _GEN_23129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23131 = 9'h97 == r_count_57_io_out ? io_r_151_b : _GEN_23130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23132 = 9'h98 == r_count_57_io_out ? io_r_152_b : _GEN_23131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23133 = 9'h99 == r_count_57_io_out ? io_r_153_b : _GEN_23132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23134 = 9'h9a == r_count_57_io_out ? io_r_154_b : _GEN_23133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23135 = 9'h9b == r_count_57_io_out ? io_r_155_b : _GEN_23134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23136 = 9'h9c == r_count_57_io_out ? io_r_156_b : _GEN_23135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23137 = 9'h9d == r_count_57_io_out ? io_r_157_b : _GEN_23136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23138 = 9'h9e == r_count_57_io_out ? io_r_158_b : _GEN_23137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23139 = 9'h9f == r_count_57_io_out ? io_r_159_b : _GEN_23138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23140 = 9'ha0 == r_count_57_io_out ? io_r_160_b : _GEN_23139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23141 = 9'ha1 == r_count_57_io_out ? io_r_161_b : _GEN_23140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23142 = 9'ha2 == r_count_57_io_out ? io_r_162_b : _GEN_23141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23143 = 9'ha3 == r_count_57_io_out ? io_r_163_b : _GEN_23142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23144 = 9'ha4 == r_count_57_io_out ? io_r_164_b : _GEN_23143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23145 = 9'ha5 == r_count_57_io_out ? io_r_165_b : _GEN_23144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23146 = 9'ha6 == r_count_57_io_out ? io_r_166_b : _GEN_23145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23147 = 9'ha7 == r_count_57_io_out ? io_r_167_b : _GEN_23146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23148 = 9'ha8 == r_count_57_io_out ? io_r_168_b : _GEN_23147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23149 = 9'ha9 == r_count_57_io_out ? io_r_169_b : _GEN_23148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23150 = 9'haa == r_count_57_io_out ? io_r_170_b : _GEN_23149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23151 = 9'hab == r_count_57_io_out ? io_r_171_b : _GEN_23150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23152 = 9'hac == r_count_57_io_out ? io_r_172_b : _GEN_23151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23153 = 9'had == r_count_57_io_out ? io_r_173_b : _GEN_23152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23154 = 9'hae == r_count_57_io_out ? io_r_174_b : _GEN_23153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23155 = 9'haf == r_count_57_io_out ? io_r_175_b : _GEN_23154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23156 = 9'hb0 == r_count_57_io_out ? io_r_176_b : _GEN_23155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23157 = 9'hb1 == r_count_57_io_out ? io_r_177_b : _GEN_23156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23158 = 9'hb2 == r_count_57_io_out ? io_r_178_b : _GEN_23157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23159 = 9'hb3 == r_count_57_io_out ? io_r_179_b : _GEN_23158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23160 = 9'hb4 == r_count_57_io_out ? io_r_180_b : _GEN_23159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23161 = 9'hb5 == r_count_57_io_out ? io_r_181_b : _GEN_23160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23162 = 9'hb6 == r_count_57_io_out ? io_r_182_b : _GEN_23161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23163 = 9'hb7 == r_count_57_io_out ? io_r_183_b : _GEN_23162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23164 = 9'hb8 == r_count_57_io_out ? io_r_184_b : _GEN_23163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23165 = 9'hb9 == r_count_57_io_out ? io_r_185_b : _GEN_23164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23166 = 9'hba == r_count_57_io_out ? io_r_186_b : _GEN_23165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23167 = 9'hbb == r_count_57_io_out ? io_r_187_b : _GEN_23166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23168 = 9'hbc == r_count_57_io_out ? io_r_188_b : _GEN_23167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23169 = 9'hbd == r_count_57_io_out ? io_r_189_b : _GEN_23168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23170 = 9'hbe == r_count_57_io_out ? io_r_190_b : _GEN_23169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23171 = 9'hbf == r_count_57_io_out ? io_r_191_b : _GEN_23170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23172 = 9'hc0 == r_count_57_io_out ? io_r_192_b : _GEN_23171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23173 = 9'hc1 == r_count_57_io_out ? io_r_193_b : _GEN_23172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23174 = 9'hc2 == r_count_57_io_out ? io_r_194_b : _GEN_23173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23175 = 9'hc3 == r_count_57_io_out ? io_r_195_b : _GEN_23174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23176 = 9'hc4 == r_count_57_io_out ? io_r_196_b : _GEN_23175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23177 = 9'hc5 == r_count_57_io_out ? io_r_197_b : _GEN_23176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23178 = 9'hc6 == r_count_57_io_out ? io_r_198_b : _GEN_23177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23179 = 9'hc7 == r_count_57_io_out ? io_r_199_b : _GEN_23178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23180 = 9'hc8 == r_count_57_io_out ? io_r_200_b : _GEN_23179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23181 = 9'hc9 == r_count_57_io_out ? io_r_201_b : _GEN_23180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23182 = 9'hca == r_count_57_io_out ? io_r_202_b : _GEN_23181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23183 = 9'hcb == r_count_57_io_out ? io_r_203_b : _GEN_23182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23184 = 9'hcc == r_count_57_io_out ? io_r_204_b : _GEN_23183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23185 = 9'hcd == r_count_57_io_out ? io_r_205_b : _GEN_23184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23186 = 9'hce == r_count_57_io_out ? io_r_206_b : _GEN_23185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23187 = 9'hcf == r_count_57_io_out ? io_r_207_b : _GEN_23186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23188 = 9'hd0 == r_count_57_io_out ? io_r_208_b : _GEN_23187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23189 = 9'hd1 == r_count_57_io_out ? io_r_209_b : _GEN_23188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23190 = 9'hd2 == r_count_57_io_out ? io_r_210_b : _GEN_23189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23191 = 9'hd3 == r_count_57_io_out ? io_r_211_b : _GEN_23190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23192 = 9'hd4 == r_count_57_io_out ? io_r_212_b : _GEN_23191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23193 = 9'hd5 == r_count_57_io_out ? io_r_213_b : _GEN_23192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23194 = 9'hd6 == r_count_57_io_out ? io_r_214_b : _GEN_23193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23195 = 9'hd7 == r_count_57_io_out ? io_r_215_b : _GEN_23194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23196 = 9'hd8 == r_count_57_io_out ? io_r_216_b : _GEN_23195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23197 = 9'hd9 == r_count_57_io_out ? io_r_217_b : _GEN_23196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23198 = 9'hda == r_count_57_io_out ? io_r_218_b : _GEN_23197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23199 = 9'hdb == r_count_57_io_out ? io_r_219_b : _GEN_23198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23200 = 9'hdc == r_count_57_io_out ? io_r_220_b : _GEN_23199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23201 = 9'hdd == r_count_57_io_out ? io_r_221_b : _GEN_23200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23202 = 9'hde == r_count_57_io_out ? io_r_222_b : _GEN_23201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23203 = 9'hdf == r_count_57_io_out ? io_r_223_b : _GEN_23202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23204 = 9'he0 == r_count_57_io_out ? io_r_224_b : _GEN_23203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23205 = 9'he1 == r_count_57_io_out ? io_r_225_b : _GEN_23204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23206 = 9'he2 == r_count_57_io_out ? io_r_226_b : _GEN_23205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23207 = 9'he3 == r_count_57_io_out ? io_r_227_b : _GEN_23206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23208 = 9'he4 == r_count_57_io_out ? io_r_228_b : _GEN_23207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23209 = 9'he5 == r_count_57_io_out ? io_r_229_b : _GEN_23208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23210 = 9'he6 == r_count_57_io_out ? io_r_230_b : _GEN_23209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23211 = 9'he7 == r_count_57_io_out ? io_r_231_b : _GEN_23210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23212 = 9'he8 == r_count_57_io_out ? io_r_232_b : _GEN_23211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23213 = 9'he9 == r_count_57_io_out ? io_r_233_b : _GEN_23212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23214 = 9'hea == r_count_57_io_out ? io_r_234_b : _GEN_23213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23215 = 9'heb == r_count_57_io_out ? io_r_235_b : _GEN_23214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23216 = 9'hec == r_count_57_io_out ? io_r_236_b : _GEN_23215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23217 = 9'hed == r_count_57_io_out ? io_r_237_b : _GEN_23216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23218 = 9'hee == r_count_57_io_out ? io_r_238_b : _GEN_23217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23219 = 9'hef == r_count_57_io_out ? io_r_239_b : _GEN_23218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23220 = 9'hf0 == r_count_57_io_out ? io_r_240_b : _GEN_23219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23221 = 9'hf1 == r_count_57_io_out ? io_r_241_b : _GEN_23220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23222 = 9'hf2 == r_count_57_io_out ? io_r_242_b : _GEN_23221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23223 = 9'hf3 == r_count_57_io_out ? io_r_243_b : _GEN_23222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23224 = 9'hf4 == r_count_57_io_out ? io_r_244_b : _GEN_23223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23225 = 9'hf5 == r_count_57_io_out ? io_r_245_b : _GEN_23224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23226 = 9'hf6 == r_count_57_io_out ? io_r_246_b : _GEN_23225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23227 = 9'hf7 == r_count_57_io_out ? io_r_247_b : _GEN_23226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23228 = 9'hf8 == r_count_57_io_out ? io_r_248_b : _GEN_23227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23229 = 9'hf9 == r_count_57_io_out ? io_r_249_b : _GEN_23228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23230 = 9'hfa == r_count_57_io_out ? io_r_250_b : _GEN_23229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23231 = 9'hfb == r_count_57_io_out ? io_r_251_b : _GEN_23230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23232 = 9'hfc == r_count_57_io_out ? io_r_252_b : _GEN_23231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23233 = 9'hfd == r_count_57_io_out ? io_r_253_b : _GEN_23232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23234 = 9'hfe == r_count_57_io_out ? io_r_254_b : _GEN_23233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23235 = 9'hff == r_count_57_io_out ? io_r_255_b : _GEN_23234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23236 = 9'h100 == r_count_57_io_out ? io_r_256_b : _GEN_23235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23237 = 9'h101 == r_count_57_io_out ? io_r_257_b : _GEN_23236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23238 = 9'h102 == r_count_57_io_out ? io_r_258_b : _GEN_23237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23239 = 9'h103 == r_count_57_io_out ? io_r_259_b : _GEN_23238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23240 = 9'h104 == r_count_57_io_out ? io_r_260_b : _GEN_23239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23241 = 9'h105 == r_count_57_io_out ? io_r_261_b : _GEN_23240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23242 = 9'h106 == r_count_57_io_out ? io_r_262_b : _GEN_23241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23243 = 9'h107 == r_count_57_io_out ? io_r_263_b : _GEN_23242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23244 = 9'h108 == r_count_57_io_out ? io_r_264_b : _GEN_23243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23245 = 9'h109 == r_count_57_io_out ? io_r_265_b : _GEN_23244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23246 = 9'h10a == r_count_57_io_out ? io_r_266_b : _GEN_23245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23247 = 9'h10b == r_count_57_io_out ? io_r_267_b : _GEN_23246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23248 = 9'h10c == r_count_57_io_out ? io_r_268_b : _GEN_23247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23249 = 9'h10d == r_count_57_io_out ? io_r_269_b : _GEN_23248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23250 = 9'h10e == r_count_57_io_out ? io_r_270_b : _GEN_23249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23251 = 9'h10f == r_count_57_io_out ? io_r_271_b : _GEN_23250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23252 = 9'h110 == r_count_57_io_out ? io_r_272_b : _GEN_23251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23253 = 9'h111 == r_count_57_io_out ? io_r_273_b : _GEN_23252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23254 = 9'h112 == r_count_57_io_out ? io_r_274_b : _GEN_23253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23255 = 9'h113 == r_count_57_io_out ? io_r_275_b : _GEN_23254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23256 = 9'h114 == r_count_57_io_out ? io_r_276_b : _GEN_23255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23257 = 9'h115 == r_count_57_io_out ? io_r_277_b : _GEN_23256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23258 = 9'h116 == r_count_57_io_out ? io_r_278_b : _GEN_23257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23259 = 9'h117 == r_count_57_io_out ? io_r_279_b : _GEN_23258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23260 = 9'h118 == r_count_57_io_out ? io_r_280_b : _GEN_23259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23261 = 9'h119 == r_count_57_io_out ? io_r_281_b : _GEN_23260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23262 = 9'h11a == r_count_57_io_out ? io_r_282_b : _GEN_23261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23263 = 9'h11b == r_count_57_io_out ? io_r_283_b : _GEN_23262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23264 = 9'h11c == r_count_57_io_out ? io_r_284_b : _GEN_23263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23265 = 9'h11d == r_count_57_io_out ? io_r_285_b : _GEN_23264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23266 = 9'h11e == r_count_57_io_out ? io_r_286_b : _GEN_23265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23267 = 9'h11f == r_count_57_io_out ? io_r_287_b : _GEN_23266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23268 = 9'h120 == r_count_57_io_out ? io_r_288_b : _GEN_23267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23269 = 9'h121 == r_count_57_io_out ? io_r_289_b : _GEN_23268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23270 = 9'h122 == r_count_57_io_out ? io_r_290_b : _GEN_23269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23271 = 9'h123 == r_count_57_io_out ? io_r_291_b : _GEN_23270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23272 = 9'h124 == r_count_57_io_out ? io_r_292_b : _GEN_23271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23273 = 9'h125 == r_count_57_io_out ? io_r_293_b : _GEN_23272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23274 = 9'h126 == r_count_57_io_out ? io_r_294_b : _GEN_23273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23275 = 9'h127 == r_count_57_io_out ? io_r_295_b : _GEN_23274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23276 = 9'h128 == r_count_57_io_out ? io_r_296_b : _GEN_23275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23277 = 9'h129 == r_count_57_io_out ? io_r_297_b : _GEN_23276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23278 = 9'h12a == r_count_57_io_out ? io_r_298_b : _GEN_23277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23279 = 9'h12b == r_count_57_io_out ? io_r_299_b : _GEN_23278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23280 = 9'h12c == r_count_57_io_out ? io_r_300_b : _GEN_23279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23281 = 9'h12d == r_count_57_io_out ? io_r_301_b : _GEN_23280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23282 = 9'h12e == r_count_57_io_out ? io_r_302_b : _GEN_23281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23283 = 9'h12f == r_count_57_io_out ? io_r_303_b : _GEN_23282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23284 = 9'h130 == r_count_57_io_out ? io_r_304_b : _GEN_23283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23285 = 9'h131 == r_count_57_io_out ? io_r_305_b : _GEN_23284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23286 = 9'h132 == r_count_57_io_out ? io_r_306_b : _GEN_23285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23287 = 9'h133 == r_count_57_io_out ? io_r_307_b : _GEN_23286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23288 = 9'h134 == r_count_57_io_out ? io_r_308_b : _GEN_23287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23289 = 9'h135 == r_count_57_io_out ? io_r_309_b : _GEN_23288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23290 = 9'h136 == r_count_57_io_out ? io_r_310_b : _GEN_23289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23291 = 9'h137 == r_count_57_io_out ? io_r_311_b : _GEN_23290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23292 = 9'h138 == r_count_57_io_out ? io_r_312_b : _GEN_23291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23293 = 9'h139 == r_count_57_io_out ? io_r_313_b : _GEN_23292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23294 = 9'h13a == r_count_57_io_out ? io_r_314_b : _GEN_23293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23295 = 9'h13b == r_count_57_io_out ? io_r_315_b : _GEN_23294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23296 = 9'h13c == r_count_57_io_out ? io_r_316_b : _GEN_23295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23297 = 9'h13d == r_count_57_io_out ? io_r_317_b : _GEN_23296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23298 = 9'h13e == r_count_57_io_out ? io_r_318_b : _GEN_23297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23299 = 9'h13f == r_count_57_io_out ? io_r_319_b : _GEN_23298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23300 = 9'h140 == r_count_57_io_out ? io_r_320_b : _GEN_23299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23301 = 9'h141 == r_count_57_io_out ? io_r_321_b : _GEN_23300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23302 = 9'h142 == r_count_57_io_out ? io_r_322_b : _GEN_23301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23303 = 9'h143 == r_count_57_io_out ? io_r_323_b : _GEN_23302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23304 = 9'h144 == r_count_57_io_out ? io_r_324_b : _GEN_23303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23305 = 9'h145 == r_count_57_io_out ? io_r_325_b : _GEN_23304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23306 = 9'h146 == r_count_57_io_out ? io_r_326_b : _GEN_23305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23307 = 9'h147 == r_count_57_io_out ? io_r_327_b : _GEN_23306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23308 = 9'h148 == r_count_57_io_out ? io_r_328_b : _GEN_23307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23309 = 9'h149 == r_count_57_io_out ? io_r_329_b : _GEN_23308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23310 = 9'h14a == r_count_57_io_out ? io_r_330_b : _GEN_23309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23311 = 9'h14b == r_count_57_io_out ? io_r_331_b : _GEN_23310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23312 = 9'h14c == r_count_57_io_out ? io_r_332_b : _GEN_23311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23313 = 9'h14d == r_count_57_io_out ? io_r_333_b : _GEN_23312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23314 = 9'h14e == r_count_57_io_out ? io_r_334_b : _GEN_23313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23315 = 9'h14f == r_count_57_io_out ? io_r_335_b : _GEN_23314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23316 = 9'h150 == r_count_57_io_out ? io_r_336_b : _GEN_23315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23317 = 9'h151 == r_count_57_io_out ? io_r_337_b : _GEN_23316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23318 = 9'h152 == r_count_57_io_out ? io_r_338_b : _GEN_23317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23319 = 9'h153 == r_count_57_io_out ? io_r_339_b : _GEN_23318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23320 = 9'h154 == r_count_57_io_out ? io_r_340_b : _GEN_23319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23321 = 9'h155 == r_count_57_io_out ? io_r_341_b : _GEN_23320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23322 = 9'h156 == r_count_57_io_out ? io_r_342_b : _GEN_23321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23323 = 9'h157 == r_count_57_io_out ? io_r_343_b : _GEN_23322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23324 = 9'h158 == r_count_57_io_out ? io_r_344_b : _GEN_23323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23325 = 9'h159 == r_count_57_io_out ? io_r_345_b : _GEN_23324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23326 = 9'h15a == r_count_57_io_out ? io_r_346_b : _GEN_23325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23327 = 9'h15b == r_count_57_io_out ? io_r_347_b : _GEN_23326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23328 = 9'h15c == r_count_57_io_out ? io_r_348_b : _GEN_23327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23329 = 9'h15d == r_count_57_io_out ? io_r_349_b : _GEN_23328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23330 = 9'h15e == r_count_57_io_out ? io_r_350_b : _GEN_23329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23331 = 9'h15f == r_count_57_io_out ? io_r_351_b : _GEN_23330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23332 = 9'h160 == r_count_57_io_out ? io_r_352_b : _GEN_23331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23333 = 9'h161 == r_count_57_io_out ? io_r_353_b : _GEN_23332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23334 = 9'h162 == r_count_57_io_out ? io_r_354_b : _GEN_23333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23335 = 9'h163 == r_count_57_io_out ? io_r_355_b : _GEN_23334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23336 = 9'h164 == r_count_57_io_out ? io_r_356_b : _GEN_23335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23337 = 9'h165 == r_count_57_io_out ? io_r_357_b : _GEN_23336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23338 = 9'h166 == r_count_57_io_out ? io_r_358_b : _GEN_23337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23339 = 9'h167 == r_count_57_io_out ? io_r_359_b : _GEN_23338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23340 = 9'h168 == r_count_57_io_out ? io_r_360_b : _GEN_23339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23341 = 9'h169 == r_count_57_io_out ? io_r_361_b : _GEN_23340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23342 = 9'h16a == r_count_57_io_out ? io_r_362_b : _GEN_23341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23343 = 9'h16b == r_count_57_io_out ? io_r_363_b : _GEN_23342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23344 = 9'h16c == r_count_57_io_out ? io_r_364_b : _GEN_23343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23345 = 9'h16d == r_count_57_io_out ? io_r_365_b : _GEN_23344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23346 = 9'h16e == r_count_57_io_out ? io_r_366_b : _GEN_23345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23347 = 9'h16f == r_count_57_io_out ? io_r_367_b : _GEN_23346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23348 = 9'h170 == r_count_57_io_out ? io_r_368_b : _GEN_23347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23349 = 9'h171 == r_count_57_io_out ? io_r_369_b : _GEN_23348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23350 = 9'h172 == r_count_57_io_out ? io_r_370_b : _GEN_23349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23351 = 9'h173 == r_count_57_io_out ? io_r_371_b : _GEN_23350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23352 = 9'h174 == r_count_57_io_out ? io_r_372_b : _GEN_23351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23353 = 9'h175 == r_count_57_io_out ? io_r_373_b : _GEN_23352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23354 = 9'h176 == r_count_57_io_out ? io_r_374_b : _GEN_23353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23355 = 9'h177 == r_count_57_io_out ? io_r_375_b : _GEN_23354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23356 = 9'h178 == r_count_57_io_out ? io_r_376_b : _GEN_23355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23357 = 9'h179 == r_count_57_io_out ? io_r_377_b : _GEN_23356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23358 = 9'h17a == r_count_57_io_out ? io_r_378_b : _GEN_23357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23359 = 9'h17b == r_count_57_io_out ? io_r_379_b : _GEN_23358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23360 = 9'h17c == r_count_57_io_out ? io_r_380_b : _GEN_23359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23361 = 9'h17d == r_count_57_io_out ? io_r_381_b : _GEN_23360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23362 = 9'h17e == r_count_57_io_out ? io_r_382_b : _GEN_23361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23363 = 9'h17f == r_count_57_io_out ? io_r_383_b : _GEN_23362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23364 = 9'h180 == r_count_57_io_out ? io_r_384_b : _GEN_23363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23365 = 9'h181 == r_count_57_io_out ? io_r_385_b : _GEN_23364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23366 = 9'h182 == r_count_57_io_out ? io_r_386_b : _GEN_23365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23367 = 9'h183 == r_count_57_io_out ? io_r_387_b : _GEN_23366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23368 = 9'h184 == r_count_57_io_out ? io_r_388_b : _GEN_23367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23369 = 9'h185 == r_count_57_io_out ? io_r_389_b : _GEN_23368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23370 = 9'h186 == r_count_57_io_out ? io_r_390_b : _GEN_23369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23371 = 9'h187 == r_count_57_io_out ? io_r_391_b : _GEN_23370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23372 = 9'h188 == r_count_57_io_out ? io_r_392_b : _GEN_23371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23373 = 9'h189 == r_count_57_io_out ? io_r_393_b : _GEN_23372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23374 = 9'h18a == r_count_57_io_out ? io_r_394_b : _GEN_23373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23375 = 9'h18b == r_count_57_io_out ? io_r_395_b : _GEN_23374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23376 = 9'h18c == r_count_57_io_out ? io_r_396_b : _GEN_23375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23377 = 9'h18d == r_count_57_io_out ? io_r_397_b : _GEN_23376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23378 = 9'h18e == r_count_57_io_out ? io_r_398_b : _GEN_23377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23381 = 9'h1 == r_count_58_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23382 = 9'h2 == r_count_58_io_out ? io_r_2_b : _GEN_23381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23383 = 9'h3 == r_count_58_io_out ? io_r_3_b : _GEN_23382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23384 = 9'h4 == r_count_58_io_out ? io_r_4_b : _GEN_23383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23385 = 9'h5 == r_count_58_io_out ? io_r_5_b : _GEN_23384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23386 = 9'h6 == r_count_58_io_out ? io_r_6_b : _GEN_23385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23387 = 9'h7 == r_count_58_io_out ? io_r_7_b : _GEN_23386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23388 = 9'h8 == r_count_58_io_out ? io_r_8_b : _GEN_23387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23389 = 9'h9 == r_count_58_io_out ? io_r_9_b : _GEN_23388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23390 = 9'ha == r_count_58_io_out ? io_r_10_b : _GEN_23389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23391 = 9'hb == r_count_58_io_out ? io_r_11_b : _GEN_23390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23392 = 9'hc == r_count_58_io_out ? io_r_12_b : _GEN_23391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23393 = 9'hd == r_count_58_io_out ? io_r_13_b : _GEN_23392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23394 = 9'he == r_count_58_io_out ? io_r_14_b : _GEN_23393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23395 = 9'hf == r_count_58_io_out ? io_r_15_b : _GEN_23394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23396 = 9'h10 == r_count_58_io_out ? io_r_16_b : _GEN_23395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23397 = 9'h11 == r_count_58_io_out ? io_r_17_b : _GEN_23396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23398 = 9'h12 == r_count_58_io_out ? io_r_18_b : _GEN_23397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23399 = 9'h13 == r_count_58_io_out ? io_r_19_b : _GEN_23398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23400 = 9'h14 == r_count_58_io_out ? io_r_20_b : _GEN_23399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23401 = 9'h15 == r_count_58_io_out ? io_r_21_b : _GEN_23400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23402 = 9'h16 == r_count_58_io_out ? io_r_22_b : _GEN_23401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23403 = 9'h17 == r_count_58_io_out ? io_r_23_b : _GEN_23402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23404 = 9'h18 == r_count_58_io_out ? io_r_24_b : _GEN_23403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23405 = 9'h19 == r_count_58_io_out ? io_r_25_b : _GEN_23404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23406 = 9'h1a == r_count_58_io_out ? io_r_26_b : _GEN_23405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23407 = 9'h1b == r_count_58_io_out ? io_r_27_b : _GEN_23406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23408 = 9'h1c == r_count_58_io_out ? io_r_28_b : _GEN_23407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23409 = 9'h1d == r_count_58_io_out ? io_r_29_b : _GEN_23408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23410 = 9'h1e == r_count_58_io_out ? io_r_30_b : _GEN_23409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23411 = 9'h1f == r_count_58_io_out ? io_r_31_b : _GEN_23410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23412 = 9'h20 == r_count_58_io_out ? io_r_32_b : _GEN_23411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23413 = 9'h21 == r_count_58_io_out ? io_r_33_b : _GEN_23412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23414 = 9'h22 == r_count_58_io_out ? io_r_34_b : _GEN_23413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23415 = 9'h23 == r_count_58_io_out ? io_r_35_b : _GEN_23414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23416 = 9'h24 == r_count_58_io_out ? io_r_36_b : _GEN_23415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23417 = 9'h25 == r_count_58_io_out ? io_r_37_b : _GEN_23416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23418 = 9'h26 == r_count_58_io_out ? io_r_38_b : _GEN_23417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23419 = 9'h27 == r_count_58_io_out ? io_r_39_b : _GEN_23418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23420 = 9'h28 == r_count_58_io_out ? io_r_40_b : _GEN_23419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23421 = 9'h29 == r_count_58_io_out ? io_r_41_b : _GEN_23420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23422 = 9'h2a == r_count_58_io_out ? io_r_42_b : _GEN_23421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23423 = 9'h2b == r_count_58_io_out ? io_r_43_b : _GEN_23422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23424 = 9'h2c == r_count_58_io_out ? io_r_44_b : _GEN_23423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23425 = 9'h2d == r_count_58_io_out ? io_r_45_b : _GEN_23424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23426 = 9'h2e == r_count_58_io_out ? io_r_46_b : _GEN_23425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23427 = 9'h2f == r_count_58_io_out ? io_r_47_b : _GEN_23426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23428 = 9'h30 == r_count_58_io_out ? io_r_48_b : _GEN_23427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23429 = 9'h31 == r_count_58_io_out ? io_r_49_b : _GEN_23428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23430 = 9'h32 == r_count_58_io_out ? io_r_50_b : _GEN_23429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23431 = 9'h33 == r_count_58_io_out ? io_r_51_b : _GEN_23430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23432 = 9'h34 == r_count_58_io_out ? io_r_52_b : _GEN_23431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23433 = 9'h35 == r_count_58_io_out ? io_r_53_b : _GEN_23432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23434 = 9'h36 == r_count_58_io_out ? io_r_54_b : _GEN_23433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23435 = 9'h37 == r_count_58_io_out ? io_r_55_b : _GEN_23434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23436 = 9'h38 == r_count_58_io_out ? io_r_56_b : _GEN_23435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23437 = 9'h39 == r_count_58_io_out ? io_r_57_b : _GEN_23436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23438 = 9'h3a == r_count_58_io_out ? io_r_58_b : _GEN_23437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23439 = 9'h3b == r_count_58_io_out ? io_r_59_b : _GEN_23438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23440 = 9'h3c == r_count_58_io_out ? io_r_60_b : _GEN_23439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23441 = 9'h3d == r_count_58_io_out ? io_r_61_b : _GEN_23440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23442 = 9'h3e == r_count_58_io_out ? io_r_62_b : _GEN_23441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23443 = 9'h3f == r_count_58_io_out ? io_r_63_b : _GEN_23442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23444 = 9'h40 == r_count_58_io_out ? io_r_64_b : _GEN_23443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23445 = 9'h41 == r_count_58_io_out ? io_r_65_b : _GEN_23444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23446 = 9'h42 == r_count_58_io_out ? io_r_66_b : _GEN_23445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23447 = 9'h43 == r_count_58_io_out ? io_r_67_b : _GEN_23446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23448 = 9'h44 == r_count_58_io_out ? io_r_68_b : _GEN_23447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23449 = 9'h45 == r_count_58_io_out ? io_r_69_b : _GEN_23448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23450 = 9'h46 == r_count_58_io_out ? io_r_70_b : _GEN_23449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23451 = 9'h47 == r_count_58_io_out ? io_r_71_b : _GEN_23450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23452 = 9'h48 == r_count_58_io_out ? io_r_72_b : _GEN_23451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23453 = 9'h49 == r_count_58_io_out ? io_r_73_b : _GEN_23452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23454 = 9'h4a == r_count_58_io_out ? io_r_74_b : _GEN_23453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23455 = 9'h4b == r_count_58_io_out ? io_r_75_b : _GEN_23454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23456 = 9'h4c == r_count_58_io_out ? io_r_76_b : _GEN_23455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23457 = 9'h4d == r_count_58_io_out ? io_r_77_b : _GEN_23456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23458 = 9'h4e == r_count_58_io_out ? io_r_78_b : _GEN_23457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23459 = 9'h4f == r_count_58_io_out ? io_r_79_b : _GEN_23458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23460 = 9'h50 == r_count_58_io_out ? io_r_80_b : _GEN_23459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23461 = 9'h51 == r_count_58_io_out ? io_r_81_b : _GEN_23460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23462 = 9'h52 == r_count_58_io_out ? io_r_82_b : _GEN_23461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23463 = 9'h53 == r_count_58_io_out ? io_r_83_b : _GEN_23462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23464 = 9'h54 == r_count_58_io_out ? io_r_84_b : _GEN_23463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23465 = 9'h55 == r_count_58_io_out ? io_r_85_b : _GEN_23464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23466 = 9'h56 == r_count_58_io_out ? io_r_86_b : _GEN_23465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23467 = 9'h57 == r_count_58_io_out ? io_r_87_b : _GEN_23466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23468 = 9'h58 == r_count_58_io_out ? io_r_88_b : _GEN_23467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23469 = 9'h59 == r_count_58_io_out ? io_r_89_b : _GEN_23468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23470 = 9'h5a == r_count_58_io_out ? io_r_90_b : _GEN_23469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23471 = 9'h5b == r_count_58_io_out ? io_r_91_b : _GEN_23470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23472 = 9'h5c == r_count_58_io_out ? io_r_92_b : _GEN_23471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23473 = 9'h5d == r_count_58_io_out ? io_r_93_b : _GEN_23472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23474 = 9'h5e == r_count_58_io_out ? io_r_94_b : _GEN_23473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23475 = 9'h5f == r_count_58_io_out ? io_r_95_b : _GEN_23474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23476 = 9'h60 == r_count_58_io_out ? io_r_96_b : _GEN_23475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23477 = 9'h61 == r_count_58_io_out ? io_r_97_b : _GEN_23476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23478 = 9'h62 == r_count_58_io_out ? io_r_98_b : _GEN_23477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23479 = 9'h63 == r_count_58_io_out ? io_r_99_b : _GEN_23478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23480 = 9'h64 == r_count_58_io_out ? io_r_100_b : _GEN_23479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23481 = 9'h65 == r_count_58_io_out ? io_r_101_b : _GEN_23480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23482 = 9'h66 == r_count_58_io_out ? io_r_102_b : _GEN_23481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23483 = 9'h67 == r_count_58_io_out ? io_r_103_b : _GEN_23482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23484 = 9'h68 == r_count_58_io_out ? io_r_104_b : _GEN_23483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23485 = 9'h69 == r_count_58_io_out ? io_r_105_b : _GEN_23484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23486 = 9'h6a == r_count_58_io_out ? io_r_106_b : _GEN_23485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23487 = 9'h6b == r_count_58_io_out ? io_r_107_b : _GEN_23486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23488 = 9'h6c == r_count_58_io_out ? io_r_108_b : _GEN_23487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23489 = 9'h6d == r_count_58_io_out ? io_r_109_b : _GEN_23488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23490 = 9'h6e == r_count_58_io_out ? io_r_110_b : _GEN_23489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23491 = 9'h6f == r_count_58_io_out ? io_r_111_b : _GEN_23490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23492 = 9'h70 == r_count_58_io_out ? io_r_112_b : _GEN_23491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23493 = 9'h71 == r_count_58_io_out ? io_r_113_b : _GEN_23492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23494 = 9'h72 == r_count_58_io_out ? io_r_114_b : _GEN_23493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23495 = 9'h73 == r_count_58_io_out ? io_r_115_b : _GEN_23494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23496 = 9'h74 == r_count_58_io_out ? io_r_116_b : _GEN_23495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23497 = 9'h75 == r_count_58_io_out ? io_r_117_b : _GEN_23496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23498 = 9'h76 == r_count_58_io_out ? io_r_118_b : _GEN_23497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23499 = 9'h77 == r_count_58_io_out ? io_r_119_b : _GEN_23498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23500 = 9'h78 == r_count_58_io_out ? io_r_120_b : _GEN_23499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23501 = 9'h79 == r_count_58_io_out ? io_r_121_b : _GEN_23500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23502 = 9'h7a == r_count_58_io_out ? io_r_122_b : _GEN_23501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23503 = 9'h7b == r_count_58_io_out ? io_r_123_b : _GEN_23502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23504 = 9'h7c == r_count_58_io_out ? io_r_124_b : _GEN_23503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23505 = 9'h7d == r_count_58_io_out ? io_r_125_b : _GEN_23504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23506 = 9'h7e == r_count_58_io_out ? io_r_126_b : _GEN_23505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23507 = 9'h7f == r_count_58_io_out ? io_r_127_b : _GEN_23506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23508 = 9'h80 == r_count_58_io_out ? io_r_128_b : _GEN_23507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23509 = 9'h81 == r_count_58_io_out ? io_r_129_b : _GEN_23508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23510 = 9'h82 == r_count_58_io_out ? io_r_130_b : _GEN_23509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23511 = 9'h83 == r_count_58_io_out ? io_r_131_b : _GEN_23510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23512 = 9'h84 == r_count_58_io_out ? io_r_132_b : _GEN_23511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23513 = 9'h85 == r_count_58_io_out ? io_r_133_b : _GEN_23512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23514 = 9'h86 == r_count_58_io_out ? io_r_134_b : _GEN_23513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23515 = 9'h87 == r_count_58_io_out ? io_r_135_b : _GEN_23514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23516 = 9'h88 == r_count_58_io_out ? io_r_136_b : _GEN_23515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23517 = 9'h89 == r_count_58_io_out ? io_r_137_b : _GEN_23516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23518 = 9'h8a == r_count_58_io_out ? io_r_138_b : _GEN_23517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23519 = 9'h8b == r_count_58_io_out ? io_r_139_b : _GEN_23518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23520 = 9'h8c == r_count_58_io_out ? io_r_140_b : _GEN_23519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23521 = 9'h8d == r_count_58_io_out ? io_r_141_b : _GEN_23520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23522 = 9'h8e == r_count_58_io_out ? io_r_142_b : _GEN_23521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23523 = 9'h8f == r_count_58_io_out ? io_r_143_b : _GEN_23522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23524 = 9'h90 == r_count_58_io_out ? io_r_144_b : _GEN_23523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23525 = 9'h91 == r_count_58_io_out ? io_r_145_b : _GEN_23524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23526 = 9'h92 == r_count_58_io_out ? io_r_146_b : _GEN_23525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23527 = 9'h93 == r_count_58_io_out ? io_r_147_b : _GEN_23526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23528 = 9'h94 == r_count_58_io_out ? io_r_148_b : _GEN_23527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23529 = 9'h95 == r_count_58_io_out ? io_r_149_b : _GEN_23528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23530 = 9'h96 == r_count_58_io_out ? io_r_150_b : _GEN_23529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23531 = 9'h97 == r_count_58_io_out ? io_r_151_b : _GEN_23530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23532 = 9'h98 == r_count_58_io_out ? io_r_152_b : _GEN_23531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23533 = 9'h99 == r_count_58_io_out ? io_r_153_b : _GEN_23532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23534 = 9'h9a == r_count_58_io_out ? io_r_154_b : _GEN_23533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23535 = 9'h9b == r_count_58_io_out ? io_r_155_b : _GEN_23534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23536 = 9'h9c == r_count_58_io_out ? io_r_156_b : _GEN_23535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23537 = 9'h9d == r_count_58_io_out ? io_r_157_b : _GEN_23536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23538 = 9'h9e == r_count_58_io_out ? io_r_158_b : _GEN_23537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23539 = 9'h9f == r_count_58_io_out ? io_r_159_b : _GEN_23538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23540 = 9'ha0 == r_count_58_io_out ? io_r_160_b : _GEN_23539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23541 = 9'ha1 == r_count_58_io_out ? io_r_161_b : _GEN_23540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23542 = 9'ha2 == r_count_58_io_out ? io_r_162_b : _GEN_23541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23543 = 9'ha3 == r_count_58_io_out ? io_r_163_b : _GEN_23542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23544 = 9'ha4 == r_count_58_io_out ? io_r_164_b : _GEN_23543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23545 = 9'ha5 == r_count_58_io_out ? io_r_165_b : _GEN_23544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23546 = 9'ha6 == r_count_58_io_out ? io_r_166_b : _GEN_23545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23547 = 9'ha7 == r_count_58_io_out ? io_r_167_b : _GEN_23546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23548 = 9'ha8 == r_count_58_io_out ? io_r_168_b : _GEN_23547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23549 = 9'ha9 == r_count_58_io_out ? io_r_169_b : _GEN_23548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23550 = 9'haa == r_count_58_io_out ? io_r_170_b : _GEN_23549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23551 = 9'hab == r_count_58_io_out ? io_r_171_b : _GEN_23550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23552 = 9'hac == r_count_58_io_out ? io_r_172_b : _GEN_23551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23553 = 9'had == r_count_58_io_out ? io_r_173_b : _GEN_23552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23554 = 9'hae == r_count_58_io_out ? io_r_174_b : _GEN_23553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23555 = 9'haf == r_count_58_io_out ? io_r_175_b : _GEN_23554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23556 = 9'hb0 == r_count_58_io_out ? io_r_176_b : _GEN_23555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23557 = 9'hb1 == r_count_58_io_out ? io_r_177_b : _GEN_23556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23558 = 9'hb2 == r_count_58_io_out ? io_r_178_b : _GEN_23557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23559 = 9'hb3 == r_count_58_io_out ? io_r_179_b : _GEN_23558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23560 = 9'hb4 == r_count_58_io_out ? io_r_180_b : _GEN_23559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23561 = 9'hb5 == r_count_58_io_out ? io_r_181_b : _GEN_23560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23562 = 9'hb6 == r_count_58_io_out ? io_r_182_b : _GEN_23561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23563 = 9'hb7 == r_count_58_io_out ? io_r_183_b : _GEN_23562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23564 = 9'hb8 == r_count_58_io_out ? io_r_184_b : _GEN_23563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23565 = 9'hb9 == r_count_58_io_out ? io_r_185_b : _GEN_23564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23566 = 9'hba == r_count_58_io_out ? io_r_186_b : _GEN_23565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23567 = 9'hbb == r_count_58_io_out ? io_r_187_b : _GEN_23566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23568 = 9'hbc == r_count_58_io_out ? io_r_188_b : _GEN_23567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23569 = 9'hbd == r_count_58_io_out ? io_r_189_b : _GEN_23568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23570 = 9'hbe == r_count_58_io_out ? io_r_190_b : _GEN_23569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23571 = 9'hbf == r_count_58_io_out ? io_r_191_b : _GEN_23570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23572 = 9'hc0 == r_count_58_io_out ? io_r_192_b : _GEN_23571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23573 = 9'hc1 == r_count_58_io_out ? io_r_193_b : _GEN_23572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23574 = 9'hc2 == r_count_58_io_out ? io_r_194_b : _GEN_23573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23575 = 9'hc3 == r_count_58_io_out ? io_r_195_b : _GEN_23574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23576 = 9'hc4 == r_count_58_io_out ? io_r_196_b : _GEN_23575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23577 = 9'hc5 == r_count_58_io_out ? io_r_197_b : _GEN_23576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23578 = 9'hc6 == r_count_58_io_out ? io_r_198_b : _GEN_23577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23579 = 9'hc7 == r_count_58_io_out ? io_r_199_b : _GEN_23578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23580 = 9'hc8 == r_count_58_io_out ? io_r_200_b : _GEN_23579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23581 = 9'hc9 == r_count_58_io_out ? io_r_201_b : _GEN_23580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23582 = 9'hca == r_count_58_io_out ? io_r_202_b : _GEN_23581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23583 = 9'hcb == r_count_58_io_out ? io_r_203_b : _GEN_23582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23584 = 9'hcc == r_count_58_io_out ? io_r_204_b : _GEN_23583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23585 = 9'hcd == r_count_58_io_out ? io_r_205_b : _GEN_23584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23586 = 9'hce == r_count_58_io_out ? io_r_206_b : _GEN_23585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23587 = 9'hcf == r_count_58_io_out ? io_r_207_b : _GEN_23586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23588 = 9'hd0 == r_count_58_io_out ? io_r_208_b : _GEN_23587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23589 = 9'hd1 == r_count_58_io_out ? io_r_209_b : _GEN_23588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23590 = 9'hd2 == r_count_58_io_out ? io_r_210_b : _GEN_23589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23591 = 9'hd3 == r_count_58_io_out ? io_r_211_b : _GEN_23590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23592 = 9'hd4 == r_count_58_io_out ? io_r_212_b : _GEN_23591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23593 = 9'hd5 == r_count_58_io_out ? io_r_213_b : _GEN_23592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23594 = 9'hd6 == r_count_58_io_out ? io_r_214_b : _GEN_23593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23595 = 9'hd7 == r_count_58_io_out ? io_r_215_b : _GEN_23594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23596 = 9'hd8 == r_count_58_io_out ? io_r_216_b : _GEN_23595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23597 = 9'hd9 == r_count_58_io_out ? io_r_217_b : _GEN_23596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23598 = 9'hda == r_count_58_io_out ? io_r_218_b : _GEN_23597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23599 = 9'hdb == r_count_58_io_out ? io_r_219_b : _GEN_23598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23600 = 9'hdc == r_count_58_io_out ? io_r_220_b : _GEN_23599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23601 = 9'hdd == r_count_58_io_out ? io_r_221_b : _GEN_23600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23602 = 9'hde == r_count_58_io_out ? io_r_222_b : _GEN_23601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23603 = 9'hdf == r_count_58_io_out ? io_r_223_b : _GEN_23602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23604 = 9'he0 == r_count_58_io_out ? io_r_224_b : _GEN_23603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23605 = 9'he1 == r_count_58_io_out ? io_r_225_b : _GEN_23604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23606 = 9'he2 == r_count_58_io_out ? io_r_226_b : _GEN_23605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23607 = 9'he3 == r_count_58_io_out ? io_r_227_b : _GEN_23606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23608 = 9'he4 == r_count_58_io_out ? io_r_228_b : _GEN_23607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23609 = 9'he5 == r_count_58_io_out ? io_r_229_b : _GEN_23608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23610 = 9'he6 == r_count_58_io_out ? io_r_230_b : _GEN_23609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23611 = 9'he7 == r_count_58_io_out ? io_r_231_b : _GEN_23610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23612 = 9'he8 == r_count_58_io_out ? io_r_232_b : _GEN_23611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23613 = 9'he9 == r_count_58_io_out ? io_r_233_b : _GEN_23612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23614 = 9'hea == r_count_58_io_out ? io_r_234_b : _GEN_23613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23615 = 9'heb == r_count_58_io_out ? io_r_235_b : _GEN_23614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23616 = 9'hec == r_count_58_io_out ? io_r_236_b : _GEN_23615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23617 = 9'hed == r_count_58_io_out ? io_r_237_b : _GEN_23616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23618 = 9'hee == r_count_58_io_out ? io_r_238_b : _GEN_23617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23619 = 9'hef == r_count_58_io_out ? io_r_239_b : _GEN_23618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23620 = 9'hf0 == r_count_58_io_out ? io_r_240_b : _GEN_23619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23621 = 9'hf1 == r_count_58_io_out ? io_r_241_b : _GEN_23620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23622 = 9'hf2 == r_count_58_io_out ? io_r_242_b : _GEN_23621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23623 = 9'hf3 == r_count_58_io_out ? io_r_243_b : _GEN_23622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23624 = 9'hf4 == r_count_58_io_out ? io_r_244_b : _GEN_23623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23625 = 9'hf5 == r_count_58_io_out ? io_r_245_b : _GEN_23624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23626 = 9'hf6 == r_count_58_io_out ? io_r_246_b : _GEN_23625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23627 = 9'hf7 == r_count_58_io_out ? io_r_247_b : _GEN_23626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23628 = 9'hf8 == r_count_58_io_out ? io_r_248_b : _GEN_23627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23629 = 9'hf9 == r_count_58_io_out ? io_r_249_b : _GEN_23628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23630 = 9'hfa == r_count_58_io_out ? io_r_250_b : _GEN_23629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23631 = 9'hfb == r_count_58_io_out ? io_r_251_b : _GEN_23630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23632 = 9'hfc == r_count_58_io_out ? io_r_252_b : _GEN_23631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23633 = 9'hfd == r_count_58_io_out ? io_r_253_b : _GEN_23632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23634 = 9'hfe == r_count_58_io_out ? io_r_254_b : _GEN_23633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23635 = 9'hff == r_count_58_io_out ? io_r_255_b : _GEN_23634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23636 = 9'h100 == r_count_58_io_out ? io_r_256_b : _GEN_23635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23637 = 9'h101 == r_count_58_io_out ? io_r_257_b : _GEN_23636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23638 = 9'h102 == r_count_58_io_out ? io_r_258_b : _GEN_23637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23639 = 9'h103 == r_count_58_io_out ? io_r_259_b : _GEN_23638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23640 = 9'h104 == r_count_58_io_out ? io_r_260_b : _GEN_23639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23641 = 9'h105 == r_count_58_io_out ? io_r_261_b : _GEN_23640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23642 = 9'h106 == r_count_58_io_out ? io_r_262_b : _GEN_23641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23643 = 9'h107 == r_count_58_io_out ? io_r_263_b : _GEN_23642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23644 = 9'h108 == r_count_58_io_out ? io_r_264_b : _GEN_23643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23645 = 9'h109 == r_count_58_io_out ? io_r_265_b : _GEN_23644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23646 = 9'h10a == r_count_58_io_out ? io_r_266_b : _GEN_23645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23647 = 9'h10b == r_count_58_io_out ? io_r_267_b : _GEN_23646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23648 = 9'h10c == r_count_58_io_out ? io_r_268_b : _GEN_23647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23649 = 9'h10d == r_count_58_io_out ? io_r_269_b : _GEN_23648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23650 = 9'h10e == r_count_58_io_out ? io_r_270_b : _GEN_23649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23651 = 9'h10f == r_count_58_io_out ? io_r_271_b : _GEN_23650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23652 = 9'h110 == r_count_58_io_out ? io_r_272_b : _GEN_23651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23653 = 9'h111 == r_count_58_io_out ? io_r_273_b : _GEN_23652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23654 = 9'h112 == r_count_58_io_out ? io_r_274_b : _GEN_23653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23655 = 9'h113 == r_count_58_io_out ? io_r_275_b : _GEN_23654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23656 = 9'h114 == r_count_58_io_out ? io_r_276_b : _GEN_23655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23657 = 9'h115 == r_count_58_io_out ? io_r_277_b : _GEN_23656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23658 = 9'h116 == r_count_58_io_out ? io_r_278_b : _GEN_23657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23659 = 9'h117 == r_count_58_io_out ? io_r_279_b : _GEN_23658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23660 = 9'h118 == r_count_58_io_out ? io_r_280_b : _GEN_23659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23661 = 9'h119 == r_count_58_io_out ? io_r_281_b : _GEN_23660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23662 = 9'h11a == r_count_58_io_out ? io_r_282_b : _GEN_23661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23663 = 9'h11b == r_count_58_io_out ? io_r_283_b : _GEN_23662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23664 = 9'h11c == r_count_58_io_out ? io_r_284_b : _GEN_23663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23665 = 9'h11d == r_count_58_io_out ? io_r_285_b : _GEN_23664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23666 = 9'h11e == r_count_58_io_out ? io_r_286_b : _GEN_23665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23667 = 9'h11f == r_count_58_io_out ? io_r_287_b : _GEN_23666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23668 = 9'h120 == r_count_58_io_out ? io_r_288_b : _GEN_23667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23669 = 9'h121 == r_count_58_io_out ? io_r_289_b : _GEN_23668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23670 = 9'h122 == r_count_58_io_out ? io_r_290_b : _GEN_23669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23671 = 9'h123 == r_count_58_io_out ? io_r_291_b : _GEN_23670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23672 = 9'h124 == r_count_58_io_out ? io_r_292_b : _GEN_23671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23673 = 9'h125 == r_count_58_io_out ? io_r_293_b : _GEN_23672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23674 = 9'h126 == r_count_58_io_out ? io_r_294_b : _GEN_23673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23675 = 9'h127 == r_count_58_io_out ? io_r_295_b : _GEN_23674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23676 = 9'h128 == r_count_58_io_out ? io_r_296_b : _GEN_23675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23677 = 9'h129 == r_count_58_io_out ? io_r_297_b : _GEN_23676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23678 = 9'h12a == r_count_58_io_out ? io_r_298_b : _GEN_23677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23679 = 9'h12b == r_count_58_io_out ? io_r_299_b : _GEN_23678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23680 = 9'h12c == r_count_58_io_out ? io_r_300_b : _GEN_23679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23681 = 9'h12d == r_count_58_io_out ? io_r_301_b : _GEN_23680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23682 = 9'h12e == r_count_58_io_out ? io_r_302_b : _GEN_23681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23683 = 9'h12f == r_count_58_io_out ? io_r_303_b : _GEN_23682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23684 = 9'h130 == r_count_58_io_out ? io_r_304_b : _GEN_23683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23685 = 9'h131 == r_count_58_io_out ? io_r_305_b : _GEN_23684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23686 = 9'h132 == r_count_58_io_out ? io_r_306_b : _GEN_23685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23687 = 9'h133 == r_count_58_io_out ? io_r_307_b : _GEN_23686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23688 = 9'h134 == r_count_58_io_out ? io_r_308_b : _GEN_23687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23689 = 9'h135 == r_count_58_io_out ? io_r_309_b : _GEN_23688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23690 = 9'h136 == r_count_58_io_out ? io_r_310_b : _GEN_23689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23691 = 9'h137 == r_count_58_io_out ? io_r_311_b : _GEN_23690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23692 = 9'h138 == r_count_58_io_out ? io_r_312_b : _GEN_23691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23693 = 9'h139 == r_count_58_io_out ? io_r_313_b : _GEN_23692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23694 = 9'h13a == r_count_58_io_out ? io_r_314_b : _GEN_23693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23695 = 9'h13b == r_count_58_io_out ? io_r_315_b : _GEN_23694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23696 = 9'h13c == r_count_58_io_out ? io_r_316_b : _GEN_23695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23697 = 9'h13d == r_count_58_io_out ? io_r_317_b : _GEN_23696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23698 = 9'h13e == r_count_58_io_out ? io_r_318_b : _GEN_23697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23699 = 9'h13f == r_count_58_io_out ? io_r_319_b : _GEN_23698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23700 = 9'h140 == r_count_58_io_out ? io_r_320_b : _GEN_23699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23701 = 9'h141 == r_count_58_io_out ? io_r_321_b : _GEN_23700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23702 = 9'h142 == r_count_58_io_out ? io_r_322_b : _GEN_23701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23703 = 9'h143 == r_count_58_io_out ? io_r_323_b : _GEN_23702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23704 = 9'h144 == r_count_58_io_out ? io_r_324_b : _GEN_23703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23705 = 9'h145 == r_count_58_io_out ? io_r_325_b : _GEN_23704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23706 = 9'h146 == r_count_58_io_out ? io_r_326_b : _GEN_23705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23707 = 9'h147 == r_count_58_io_out ? io_r_327_b : _GEN_23706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23708 = 9'h148 == r_count_58_io_out ? io_r_328_b : _GEN_23707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23709 = 9'h149 == r_count_58_io_out ? io_r_329_b : _GEN_23708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23710 = 9'h14a == r_count_58_io_out ? io_r_330_b : _GEN_23709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23711 = 9'h14b == r_count_58_io_out ? io_r_331_b : _GEN_23710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23712 = 9'h14c == r_count_58_io_out ? io_r_332_b : _GEN_23711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23713 = 9'h14d == r_count_58_io_out ? io_r_333_b : _GEN_23712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23714 = 9'h14e == r_count_58_io_out ? io_r_334_b : _GEN_23713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23715 = 9'h14f == r_count_58_io_out ? io_r_335_b : _GEN_23714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23716 = 9'h150 == r_count_58_io_out ? io_r_336_b : _GEN_23715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23717 = 9'h151 == r_count_58_io_out ? io_r_337_b : _GEN_23716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23718 = 9'h152 == r_count_58_io_out ? io_r_338_b : _GEN_23717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23719 = 9'h153 == r_count_58_io_out ? io_r_339_b : _GEN_23718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23720 = 9'h154 == r_count_58_io_out ? io_r_340_b : _GEN_23719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23721 = 9'h155 == r_count_58_io_out ? io_r_341_b : _GEN_23720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23722 = 9'h156 == r_count_58_io_out ? io_r_342_b : _GEN_23721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23723 = 9'h157 == r_count_58_io_out ? io_r_343_b : _GEN_23722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23724 = 9'h158 == r_count_58_io_out ? io_r_344_b : _GEN_23723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23725 = 9'h159 == r_count_58_io_out ? io_r_345_b : _GEN_23724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23726 = 9'h15a == r_count_58_io_out ? io_r_346_b : _GEN_23725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23727 = 9'h15b == r_count_58_io_out ? io_r_347_b : _GEN_23726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23728 = 9'h15c == r_count_58_io_out ? io_r_348_b : _GEN_23727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23729 = 9'h15d == r_count_58_io_out ? io_r_349_b : _GEN_23728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23730 = 9'h15e == r_count_58_io_out ? io_r_350_b : _GEN_23729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23731 = 9'h15f == r_count_58_io_out ? io_r_351_b : _GEN_23730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23732 = 9'h160 == r_count_58_io_out ? io_r_352_b : _GEN_23731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23733 = 9'h161 == r_count_58_io_out ? io_r_353_b : _GEN_23732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23734 = 9'h162 == r_count_58_io_out ? io_r_354_b : _GEN_23733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23735 = 9'h163 == r_count_58_io_out ? io_r_355_b : _GEN_23734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23736 = 9'h164 == r_count_58_io_out ? io_r_356_b : _GEN_23735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23737 = 9'h165 == r_count_58_io_out ? io_r_357_b : _GEN_23736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23738 = 9'h166 == r_count_58_io_out ? io_r_358_b : _GEN_23737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23739 = 9'h167 == r_count_58_io_out ? io_r_359_b : _GEN_23738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23740 = 9'h168 == r_count_58_io_out ? io_r_360_b : _GEN_23739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23741 = 9'h169 == r_count_58_io_out ? io_r_361_b : _GEN_23740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23742 = 9'h16a == r_count_58_io_out ? io_r_362_b : _GEN_23741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23743 = 9'h16b == r_count_58_io_out ? io_r_363_b : _GEN_23742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23744 = 9'h16c == r_count_58_io_out ? io_r_364_b : _GEN_23743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23745 = 9'h16d == r_count_58_io_out ? io_r_365_b : _GEN_23744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23746 = 9'h16e == r_count_58_io_out ? io_r_366_b : _GEN_23745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23747 = 9'h16f == r_count_58_io_out ? io_r_367_b : _GEN_23746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23748 = 9'h170 == r_count_58_io_out ? io_r_368_b : _GEN_23747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23749 = 9'h171 == r_count_58_io_out ? io_r_369_b : _GEN_23748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23750 = 9'h172 == r_count_58_io_out ? io_r_370_b : _GEN_23749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23751 = 9'h173 == r_count_58_io_out ? io_r_371_b : _GEN_23750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23752 = 9'h174 == r_count_58_io_out ? io_r_372_b : _GEN_23751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23753 = 9'h175 == r_count_58_io_out ? io_r_373_b : _GEN_23752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23754 = 9'h176 == r_count_58_io_out ? io_r_374_b : _GEN_23753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23755 = 9'h177 == r_count_58_io_out ? io_r_375_b : _GEN_23754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23756 = 9'h178 == r_count_58_io_out ? io_r_376_b : _GEN_23755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23757 = 9'h179 == r_count_58_io_out ? io_r_377_b : _GEN_23756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23758 = 9'h17a == r_count_58_io_out ? io_r_378_b : _GEN_23757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23759 = 9'h17b == r_count_58_io_out ? io_r_379_b : _GEN_23758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23760 = 9'h17c == r_count_58_io_out ? io_r_380_b : _GEN_23759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23761 = 9'h17d == r_count_58_io_out ? io_r_381_b : _GEN_23760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23762 = 9'h17e == r_count_58_io_out ? io_r_382_b : _GEN_23761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23763 = 9'h17f == r_count_58_io_out ? io_r_383_b : _GEN_23762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23764 = 9'h180 == r_count_58_io_out ? io_r_384_b : _GEN_23763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23765 = 9'h181 == r_count_58_io_out ? io_r_385_b : _GEN_23764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23766 = 9'h182 == r_count_58_io_out ? io_r_386_b : _GEN_23765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23767 = 9'h183 == r_count_58_io_out ? io_r_387_b : _GEN_23766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23768 = 9'h184 == r_count_58_io_out ? io_r_388_b : _GEN_23767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23769 = 9'h185 == r_count_58_io_out ? io_r_389_b : _GEN_23768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23770 = 9'h186 == r_count_58_io_out ? io_r_390_b : _GEN_23769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23771 = 9'h187 == r_count_58_io_out ? io_r_391_b : _GEN_23770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23772 = 9'h188 == r_count_58_io_out ? io_r_392_b : _GEN_23771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23773 = 9'h189 == r_count_58_io_out ? io_r_393_b : _GEN_23772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23774 = 9'h18a == r_count_58_io_out ? io_r_394_b : _GEN_23773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23775 = 9'h18b == r_count_58_io_out ? io_r_395_b : _GEN_23774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23776 = 9'h18c == r_count_58_io_out ? io_r_396_b : _GEN_23775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23777 = 9'h18d == r_count_58_io_out ? io_r_397_b : _GEN_23776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23778 = 9'h18e == r_count_58_io_out ? io_r_398_b : _GEN_23777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23781 = 9'h1 == r_count_59_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23782 = 9'h2 == r_count_59_io_out ? io_r_2_b : _GEN_23781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23783 = 9'h3 == r_count_59_io_out ? io_r_3_b : _GEN_23782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23784 = 9'h4 == r_count_59_io_out ? io_r_4_b : _GEN_23783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23785 = 9'h5 == r_count_59_io_out ? io_r_5_b : _GEN_23784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23786 = 9'h6 == r_count_59_io_out ? io_r_6_b : _GEN_23785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23787 = 9'h7 == r_count_59_io_out ? io_r_7_b : _GEN_23786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23788 = 9'h8 == r_count_59_io_out ? io_r_8_b : _GEN_23787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23789 = 9'h9 == r_count_59_io_out ? io_r_9_b : _GEN_23788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23790 = 9'ha == r_count_59_io_out ? io_r_10_b : _GEN_23789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23791 = 9'hb == r_count_59_io_out ? io_r_11_b : _GEN_23790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23792 = 9'hc == r_count_59_io_out ? io_r_12_b : _GEN_23791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23793 = 9'hd == r_count_59_io_out ? io_r_13_b : _GEN_23792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23794 = 9'he == r_count_59_io_out ? io_r_14_b : _GEN_23793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23795 = 9'hf == r_count_59_io_out ? io_r_15_b : _GEN_23794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23796 = 9'h10 == r_count_59_io_out ? io_r_16_b : _GEN_23795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23797 = 9'h11 == r_count_59_io_out ? io_r_17_b : _GEN_23796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23798 = 9'h12 == r_count_59_io_out ? io_r_18_b : _GEN_23797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23799 = 9'h13 == r_count_59_io_out ? io_r_19_b : _GEN_23798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23800 = 9'h14 == r_count_59_io_out ? io_r_20_b : _GEN_23799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23801 = 9'h15 == r_count_59_io_out ? io_r_21_b : _GEN_23800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23802 = 9'h16 == r_count_59_io_out ? io_r_22_b : _GEN_23801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23803 = 9'h17 == r_count_59_io_out ? io_r_23_b : _GEN_23802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23804 = 9'h18 == r_count_59_io_out ? io_r_24_b : _GEN_23803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23805 = 9'h19 == r_count_59_io_out ? io_r_25_b : _GEN_23804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23806 = 9'h1a == r_count_59_io_out ? io_r_26_b : _GEN_23805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23807 = 9'h1b == r_count_59_io_out ? io_r_27_b : _GEN_23806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23808 = 9'h1c == r_count_59_io_out ? io_r_28_b : _GEN_23807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23809 = 9'h1d == r_count_59_io_out ? io_r_29_b : _GEN_23808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23810 = 9'h1e == r_count_59_io_out ? io_r_30_b : _GEN_23809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23811 = 9'h1f == r_count_59_io_out ? io_r_31_b : _GEN_23810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23812 = 9'h20 == r_count_59_io_out ? io_r_32_b : _GEN_23811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23813 = 9'h21 == r_count_59_io_out ? io_r_33_b : _GEN_23812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23814 = 9'h22 == r_count_59_io_out ? io_r_34_b : _GEN_23813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23815 = 9'h23 == r_count_59_io_out ? io_r_35_b : _GEN_23814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23816 = 9'h24 == r_count_59_io_out ? io_r_36_b : _GEN_23815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23817 = 9'h25 == r_count_59_io_out ? io_r_37_b : _GEN_23816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23818 = 9'h26 == r_count_59_io_out ? io_r_38_b : _GEN_23817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23819 = 9'h27 == r_count_59_io_out ? io_r_39_b : _GEN_23818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23820 = 9'h28 == r_count_59_io_out ? io_r_40_b : _GEN_23819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23821 = 9'h29 == r_count_59_io_out ? io_r_41_b : _GEN_23820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23822 = 9'h2a == r_count_59_io_out ? io_r_42_b : _GEN_23821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23823 = 9'h2b == r_count_59_io_out ? io_r_43_b : _GEN_23822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23824 = 9'h2c == r_count_59_io_out ? io_r_44_b : _GEN_23823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23825 = 9'h2d == r_count_59_io_out ? io_r_45_b : _GEN_23824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23826 = 9'h2e == r_count_59_io_out ? io_r_46_b : _GEN_23825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23827 = 9'h2f == r_count_59_io_out ? io_r_47_b : _GEN_23826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23828 = 9'h30 == r_count_59_io_out ? io_r_48_b : _GEN_23827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23829 = 9'h31 == r_count_59_io_out ? io_r_49_b : _GEN_23828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23830 = 9'h32 == r_count_59_io_out ? io_r_50_b : _GEN_23829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23831 = 9'h33 == r_count_59_io_out ? io_r_51_b : _GEN_23830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23832 = 9'h34 == r_count_59_io_out ? io_r_52_b : _GEN_23831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23833 = 9'h35 == r_count_59_io_out ? io_r_53_b : _GEN_23832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23834 = 9'h36 == r_count_59_io_out ? io_r_54_b : _GEN_23833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23835 = 9'h37 == r_count_59_io_out ? io_r_55_b : _GEN_23834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23836 = 9'h38 == r_count_59_io_out ? io_r_56_b : _GEN_23835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23837 = 9'h39 == r_count_59_io_out ? io_r_57_b : _GEN_23836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23838 = 9'h3a == r_count_59_io_out ? io_r_58_b : _GEN_23837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23839 = 9'h3b == r_count_59_io_out ? io_r_59_b : _GEN_23838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23840 = 9'h3c == r_count_59_io_out ? io_r_60_b : _GEN_23839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23841 = 9'h3d == r_count_59_io_out ? io_r_61_b : _GEN_23840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23842 = 9'h3e == r_count_59_io_out ? io_r_62_b : _GEN_23841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23843 = 9'h3f == r_count_59_io_out ? io_r_63_b : _GEN_23842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23844 = 9'h40 == r_count_59_io_out ? io_r_64_b : _GEN_23843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23845 = 9'h41 == r_count_59_io_out ? io_r_65_b : _GEN_23844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23846 = 9'h42 == r_count_59_io_out ? io_r_66_b : _GEN_23845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23847 = 9'h43 == r_count_59_io_out ? io_r_67_b : _GEN_23846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23848 = 9'h44 == r_count_59_io_out ? io_r_68_b : _GEN_23847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23849 = 9'h45 == r_count_59_io_out ? io_r_69_b : _GEN_23848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23850 = 9'h46 == r_count_59_io_out ? io_r_70_b : _GEN_23849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23851 = 9'h47 == r_count_59_io_out ? io_r_71_b : _GEN_23850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23852 = 9'h48 == r_count_59_io_out ? io_r_72_b : _GEN_23851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23853 = 9'h49 == r_count_59_io_out ? io_r_73_b : _GEN_23852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23854 = 9'h4a == r_count_59_io_out ? io_r_74_b : _GEN_23853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23855 = 9'h4b == r_count_59_io_out ? io_r_75_b : _GEN_23854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23856 = 9'h4c == r_count_59_io_out ? io_r_76_b : _GEN_23855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23857 = 9'h4d == r_count_59_io_out ? io_r_77_b : _GEN_23856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23858 = 9'h4e == r_count_59_io_out ? io_r_78_b : _GEN_23857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23859 = 9'h4f == r_count_59_io_out ? io_r_79_b : _GEN_23858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23860 = 9'h50 == r_count_59_io_out ? io_r_80_b : _GEN_23859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23861 = 9'h51 == r_count_59_io_out ? io_r_81_b : _GEN_23860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23862 = 9'h52 == r_count_59_io_out ? io_r_82_b : _GEN_23861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23863 = 9'h53 == r_count_59_io_out ? io_r_83_b : _GEN_23862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23864 = 9'h54 == r_count_59_io_out ? io_r_84_b : _GEN_23863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23865 = 9'h55 == r_count_59_io_out ? io_r_85_b : _GEN_23864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23866 = 9'h56 == r_count_59_io_out ? io_r_86_b : _GEN_23865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23867 = 9'h57 == r_count_59_io_out ? io_r_87_b : _GEN_23866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23868 = 9'h58 == r_count_59_io_out ? io_r_88_b : _GEN_23867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23869 = 9'h59 == r_count_59_io_out ? io_r_89_b : _GEN_23868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23870 = 9'h5a == r_count_59_io_out ? io_r_90_b : _GEN_23869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23871 = 9'h5b == r_count_59_io_out ? io_r_91_b : _GEN_23870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23872 = 9'h5c == r_count_59_io_out ? io_r_92_b : _GEN_23871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23873 = 9'h5d == r_count_59_io_out ? io_r_93_b : _GEN_23872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23874 = 9'h5e == r_count_59_io_out ? io_r_94_b : _GEN_23873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23875 = 9'h5f == r_count_59_io_out ? io_r_95_b : _GEN_23874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23876 = 9'h60 == r_count_59_io_out ? io_r_96_b : _GEN_23875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23877 = 9'h61 == r_count_59_io_out ? io_r_97_b : _GEN_23876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23878 = 9'h62 == r_count_59_io_out ? io_r_98_b : _GEN_23877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23879 = 9'h63 == r_count_59_io_out ? io_r_99_b : _GEN_23878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23880 = 9'h64 == r_count_59_io_out ? io_r_100_b : _GEN_23879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23881 = 9'h65 == r_count_59_io_out ? io_r_101_b : _GEN_23880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23882 = 9'h66 == r_count_59_io_out ? io_r_102_b : _GEN_23881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23883 = 9'h67 == r_count_59_io_out ? io_r_103_b : _GEN_23882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23884 = 9'h68 == r_count_59_io_out ? io_r_104_b : _GEN_23883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23885 = 9'h69 == r_count_59_io_out ? io_r_105_b : _GEN_23884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23886 = 9'h6a == r_count_59_io_out ? io_r_106_b : _GEN_23885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23887 = 9'h6b == r_count_59_io_out ? io_r_107_b : _GEN_23886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23888 = 9'h6c == r_count_59_io_out ? io_r_108_b : _GEN_23887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23889 = 9'h6d == r_count_59_io_out ? io_r_109_b : _GEN_23888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23890 = 9'h6e == r_count_59_io_out ? io_r_110_b : _GEN_23889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23891 = 9'h6f == r_count_59_io_out ? io_r_111_b : _GEN_23890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23892 = 9'h70 == r_count_59_io_out ? io_r_112_b : _GEN_23891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23893 = 9'h71 == r_count_59_io_out ? io_r_113_b : _GEN_23892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23894 = 9'h72 == r_count_59_io_out ? io_r_114_b : _GEN_23893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23895 = 9'h73 == r_count_59_io_out ? io_r_115_b : _GEN_23894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23896 = 9'h74 == r_count_59_io_out ? io_r_116_b : _GEN_23895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23897 = 9'h75 == r_count_59_io_out ? io_r_117_b : _GEN_23896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23898 = 9'h76 == r_count_59_io_out ? io_r_118_b : _GEN_23897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23899 = 9'h77 == r_count_59_io_out ? io_r_119_b : _GEN_23898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23900 = 9'h78 == r_count_59_io_out ? io_r_120_b : _GEN_23899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23901 = 9'h79 == r_count_59_io_out ? io_r_121_b : _GEN_23900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23902 = 9'h7a == r_count_59_io_out ? io_r_122_b : _GEN_23901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23903 = 9'h7b == r_count_59_io_out ? io_r_123_b : _GEN_23902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23904 = 9'h7c == r_count_59_io_out ? io_r_124_b : _GEN_23903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23905 = 9'h7d == r_count_59_io_out ? io_r_125_b : _GEN_23904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23906 = 9'h7e == r_count_59_io_out ? io_r_126_b : _GEN_23905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23907 = 9'h7f == r_count_59_io_out ? io_r_127_b : _GEN_23906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23908 = 9'h80 == r_count_59_io_out ? io_r_128_b : _GEN_23907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23909 = 9'h81 == r_count_59_io_out ? io_r_129_b : _GEN_23908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23910 = 9'h82 == r_count_59_io_out ? io_r_130_b : _GEN_23909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23911 = 9'h83 == r_count_59_io_out ? io_r_131_b : _GEN_23910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23912 = 9'h84 == r_count_59_io_out ? io_r_132_b : _GEN_23911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23913 = 9'h85 == r_count_59_io_out ? io_r_133_b : _GEN_23912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23914 = 9'h86 == r_count_59_io_out ? io_r_134_b : _GEN_23913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23915 = 9'h87 == r_count_59_io_out ? io_r_135_b : _GEN_23914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23916 = 9'h88 == r_count_59_io_out ? io_r_136_b : _GEN_23915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23917 = 9'h89 == r_count_59_io_out ? io_r_137_b : _GEN_23916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23918 = 9'h8a == r_count_59_io_out ? io_r_138_b : _GEN_23917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23919 = 9'h8b == r_count_59_io_out ? io_r_139_b : _GEN_23918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23920 = 9'h8c == r_count_59_io_out ? io_r_140_b : _GEN_23919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23921 = 9'h8d == r_count_59_io_out ? io_r_141_b : _GEN_23920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23922 = 9'h8e == r_count_59_io_out ? io_r_142_b : _GEN_23921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23923 = 9'h8f == r_count_59_io_out ? io_r_143_b : _GEN_23922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23924 = 9'h90 == r_count_59_io_out ? io_r_144_b : _GEN_23923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23925 = 9'h91 == r_count_59_io_out ? io_r_145_b : _GEN_23924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23926 = 9'h92 == r_count_59_io_out ? io_r_146_b : _GEN_23925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23927 = 9'h93 == r_count_59_io_out ? io_r_147_b : _GEN_23926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23928 = 9'h94 == r_count_59_io_out ? io_r_148_b : _GEN_23927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23929 = 9'h95 == r_count_59_io_out ? io_r_149_b : _GEN_23928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23930 = 9'h96 == r_count_59_io_out ? io_r_150_b : _GEN_23929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23931 = 9'h97 == r_count_59_io_out ? io_r_151_b : _GEN_23930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23932 = 9'h98 == r_count_59_io_out ? io_r_152_b : _GEN_23931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23933 = 9'h99 == r_count_59_io_out ? io_r_153_b : _GEN_23932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23934 = 9'h9a == r_count_59_io_out ? io_r_154_b : _GEN_23933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23935 = 9'h9b == r_count_59_io_out ? io_r_155_b : _GEN_23934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23936 = 9'h9c == r_count_59_io_out ? io_r_156_b : _GEN_23935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23937 = 9'h9d == r_count_59_io_out ? io_r_157_b : _GEN_23936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23938 = 9'h9e == r_count_59_io_out ? io_r_158_b : _GEN_23937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23939 = 9'h9f == r_count_59_io_out ? io_r_159_b : _GEN_23938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23940 = 9'ha0 == r_count_59_io_out ? io_r_160_b : _GEN_23939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23941 = 9'ha1 == r_count_59_io_out ? io_r_161_b : _GEN_23940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23942 = 9'ha2 == r_count_59_io_out ? io_r_162_b : _GEN_23941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23943 = 9'ha3 == r_count_59_io_out ? io_r_163_b : _GEN_23942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23944 = 9'ha4 == r_count_59_io_out ? io_r_164_b : _GEN_23943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23945 = 9'ha5 == r_count_59_io_out ? io_r_165_b : _GEN_23944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23946 = 9'ha6 == r_count_59_io_out ? io_r_166_b : _GEN_23945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23947 = 9'ha7 == r_count_59_io_out ? io_r_167_b : _GEN_23946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23948 = 9'ha8 == r_count_59_io_out ? io_r_168_b : _GEN_23947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23949 = 9'ha9 == r_count_59_io_out ? io_r_169_b : _GEN_23948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23950 = 9'haa == r_count_59_io_out ? io_r_170_b : _GEN_23949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23951 = 9'hab == r_count_59_io_out ? io_r_171_b : _GEN_23950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23952 = 9'hac == r_count_59_io_out ? io_r_172_b : _GEN_23951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23953 = 9'had == r_count_59_io_out ? io_r_173_b : _GEN_23952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23954 = 9'hae == r_count_59_io_out ? io_r_174_b : _GEN_23953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23955 = 9'haf == r_count_59_io_out ? io_r_175_b : _GEN_23954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23956 = 9'hb0 == r_count_59_io_out ? io_r_176_b : _GEN_23955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23957 = 9'hb1 == r_count_59_io_out ? io_r_177_b : _GEN_23956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23958 = 9'hb2 == r_count_59_io_out ? io_r_178_b : _GEN_23957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23959 = 9'hb3 == r_count_59_io_out ? io_r_179_b : _GEN_23958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23960 = 9'hb4 == r_count_59_io_out ? io_r_180_b : _GEN_23959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23961 = 9'hb5 == r_count_59_io_out ? io_r_181_b : _GEN_23960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23962 = 9'hb6 == r_count_59_io_out ? io_r_182_b : _GEN_23961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23963 = 9'hb7 == r_count_59_io_out ? io_r_183_b : _GEN_23962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23964 = 9'hb8 == r_count_59_io_out ? io_r_184_b : _GEN_23963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23965 = 9'hb9 == r_count_59_io_out ? io_r_185_b : _GEN_23964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23966 = 9'hba == r_count_59_io_out ? io_r_186_b : _GEN_23965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23967 = 9'hbb == r_count_59_io_out ? io_r_187_b : _GEN_23966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23968 = 9'hbc == r_count_59_io_out ? io_r_188_b : _GEN_23967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23969 = 9'hbd == r_count_59_io_out ? io_r_189_b : _GEN_23968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23970 = 9'hbe == r_count_59_io_out ? io_r_190_b : _GEN_23969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23971 = 9'hbf == r_count_59_io_out ? io_r_191_b : _GEN_23970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23972 = 9'hc0 == r_count_59_io_out ? io_r_192_b : _GEN_23971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23973 = 9'hc1 == r_count_59_io_out ? io_r_193_b : _GEN_23972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23974 = 9'hc2 == r_count_59_io_out ? io_r_194_b : _GEN_23973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23975 = 9'hc3 == r_count_59_io_out ? io_r_195_b : _GEN_23974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23976 = 9'hc4 == r_count_59_io_out ? io_r_196_b : _GEN_23975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23977 = 9'hc5 == r_count_59_io_out ? io_r_197_b : _GEN_23976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23978 = 9'hc6 == r_count_59_io_out ? io_r_198_b : _GEN_23977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23979 = 9'hc7 == r_count_59_io_out ? io_r_199_b : _GEN_23978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23980 = 9'hc8 == r_count_59_io_out ? io_r_200_b : _GEN_23979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23981 = 9'hc9 == r_count_59_io_out ? io_r_201_b : _GEN_23980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23982 = 9'hca == r_count_59_io_out ? io_r_202_b : _GEN_23981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23983 = 9'hcb == r_count_59_io_out ? io_r_203_b : _GEN_23982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23984 = 9'hcc == r_count_59_io_out ? io_r_204_b : _GEN_23983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23985 = 9'hcd == r_count_59_io_out ? io_r_205_b : _GEN_23984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23986 = 9'hce == r_count_59_io_out ? io_r_206_b : _GEN_23985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23987 = 9'hcf == r_count_59_io_out ? io_r_207_b : _GEN_23986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23988 = 9'hd0 == r_count_59_io_out ? io_r_208_b : _GEN_23987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23989 = 9'hd1 == r_count_59_io_out ? io_r_209_b : _GEN_23988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23990 = 9'hd2 == r_count_59_io_out ? io_r_210_b : _GEN_23989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23991 = 9'hd3 == r_count_59_io_out ? io_r_211_b : _GEN_23990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23992 = 9'hd4 == r_count_59_io_out ? io_r_212_b : _GEN_23991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23993 = 9'hd5 == r_count_59_io_out ? io_r_213_b : _GEN_23992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23994 = 9'hd6 == r_count_59_io_out ? io_r_214_b : _GEN_23993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23995 = 9'hd7 == r_count_59_io_out ? io_r_215_b : _GEN_23994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23996 = 9'hd8 == r_count_59_io_out ? io_r_216_b : _GEN_23995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23997 = 9'hd9 == r_count_59_io_out ? io_r_217_b : _GEN_23996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23998 = 9'hda == r_count_59_io_out ? io_r_218_b : _GEN_23997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_23999 = 9'hdb == r_count_59_io_out ? io_r_219_b : _GEN_23998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24000 = 9'hdc == r_count_59_io_out ? io_r_220_b : _GEN_23999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24001 = 9'hdd == r_count_59_io_out ? io_r_221_b : _GEN_24000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24002 = 9'hde == r_count_59_io_out ? io_r_222_b : _GEN_24001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24003 = 9'hdf == r_count_59_io_out ? io_r_223_b : _GEN_24002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24004 = 9'he0 == r_count_59_io_out ? io_r_224_b : _GEN_24003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24005 = 9'he1 == r_count_59_io_out ? io_r_225_b : _GEN_24004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24006 = 9'he2 == r_count_59_io_out ? io_r_226_b : _GEN_24005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24007 = 9'he3 == r_count_59_io_out ? io_r_227_b : _GEN_24006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24008 = 9'he4 == r_count_59_io_out ? io_r_228_b : _GEN_24007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24009 = 9'he5 == r_count_59_io_out ? io_r_229_b : _GEN_24008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24010 = 9'he6 == r_count_59_io_out ? io_r_230_b : _GEN_24009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24011 = 9'he7 == r_count_59_io_out ? io_r_231_b : _GEN_24010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24012 = 9'he8 == r_count_59_io_out ? io_r_232_b : _GEN_24011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24013 = 9'he9 == r_count_59_io_out ? io_r_233_b : _GEN_24012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24014 = 9'hea == r_count_59_io_out ? io_r_234_b : _GEN_24013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24015 = 9'heb == r_count_59_io_out ? io_r_235_b : _GEN_24014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24016 = 9'hec == r_count_59_io_out ? io_r_236_b : _GEN_24015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24017 = 9'hed == r_count_59_io_out ? io_r_237_b : _GEN_24016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24018 = 9'hee == r_count_59_io_out ? io_r_238_b : _GEN_24017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24019 = 9'hef == r_count_59_io_out ? io_r_239_b : _GEN_24018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24020 = 9'hf0 == r_count_59_io_out ? io_r_240_b : _GEN_24019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24021 = 9'hf1 == r_count_59_io_out ? io_r_241_b : _GEN_24020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24022 = 9'hf2 == r_count_59_io_out ? io_r_242_b : _GEN_24021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24023 = 9'hf3 == r_count_59_io_out ? io_r_243_b : _GEN_24022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24024 = 9'hf4 == r_count_59_io_out ? io_r_244_b : _GEN_24023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24025 = 9'hf5 == r_count_59_io_out ? io_r_245_b : _GEN_24024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24026 = 9'hf6 == r_count_59_io_out ? io_r_246_b : _GEN_24025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24027 = 9'hf7 == r_count_59_io_out ? io_r_247_b : _GEN_24026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24028 = 9'hf8 == r_count_59_io_out ? io_r_248_b : _GEN_24027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24029 = 9'hf9 == r_count_59_io_out ? io_r_249_b : _GEN_24028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24030 = 9'hfa == r_count_59_io_out ? io_r_250_b : _GEN_24029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24031 = 9'hfb == r_count_59_io_out ? io_r_251_b : _GEN_24030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24032 = 9'hfc == r_count_59_io_out ? io_r_252_b : _GEN_24031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24033 = 9'hfd == r_count_59_io_out ? io_r_253_b : _GEN_24032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24034 = 9'hfe == r_count_59_io_out ? io_r_254_b : _GEN_24033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24035 = 9'hff == r_count_59_io_out ? io_r_255_b : _GEN_24034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24036 = 9'h100 == r_count_59_io_out ? io_r_256_b : _GEN_24035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24037 = 9'h101 == r_count_59_io_out ? io_r_257_b : _GEN_24036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24038 = 9'h102 == r_count_59_io_out ? io_r_258_b : _GEN_24037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24039 = 9'h103 == r_count_59_io_out ? io_r_259_b : _GEN_24038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24040 = 9'h104 == r_count_59_io_out ? io_r_260_b : _GEN_24039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24041 = 9'h105 == r_count_59_io_out ? io_r_261_b : _GEN_24040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24042 = 9'h106 == r_count_59_io_out ? io_r_262_b : _GEN_24041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24043 = 9'h107 == r_count_59_io_out ? io_r_263_b : _GEN_24042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24044 = 9'h108 == r_count_59_io_out ? io_r_264_b : _GEN_24043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24045 = 9'h109 == r_count_59_io_out ? io_r_265_b : _GEN_24044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24046 = 9'h10a == r_count_59_io_out ? io_r_266_b : _GEN_24045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24047 = 9'h10b == r_count_59_io_out ? io_r_267_b : _GEN_24046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24048 = 9'h10c == r_count_59_io_out ? io_r_268_b : _GEN_24047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24049 = 9'h10d == r_count_59_io_out ? io_r_269_b : _GEN_24048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24050 = 9'h10e == r_count_59_io_out ? io_r_270_b : _GEN_24049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24051 = 9'h10f == r_count_59_io_out ? io_r_271_b : _GEN_24050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24052 = 9'h110 == r_count_59_io_out ? io_r_272_b : _GEN_24051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24053 = 9'h111 == r_count_59_io_out ? io_r_273_b : _GEN_24052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24054 = 9'h112 == r_count_59_io_out ? io_r_274_b : _GEN_24053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24055 = 9'h113 == r_count_59_io_out ? io_r_275_b : _GEN_24054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24056 = 9'h114 == r_count_59_io_out ? io_r_276_b : _GEN_24055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24057 = 9'h115 == r_count_59_io_out ? io_r_277_b : _GEN_24056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24058 = 9'h116 == r_count_59_io_out ? io_r_278_b : _GEN_24057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24059 = 9'h117 == r_count_59_io_out ? io_r_279_b : _GEN_24058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24060 = 9'h118 == r_count_59_io_out ? io_r_280_b : _GEN_24059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24061 = 9'h119 == r_count_59_io_out ? io_r_281_b : _GEN_24060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24062 = 9'h11a == r_count_59_io_out ? io_r_282_b : _GEN_24061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24063 = 9'h11b == r_count_59_io_out ? io_r_283_b : _GEN_24062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24064 = 9'h11c == r_count_59_io_out ? io_r_284_b : _GEN_24063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24065 = 9'h11d == r_count_59_io_out ? io_r_285_b : _GEN_24064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24066 = 9'h11e == r_count_59_io_out ? io_r_286_b : _GEN_24065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24067 = 9'h11f == r_count_59_io_out ? io_r_287_b : _GEN_24066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24068 = 9'h120 == r_count_59_io_out ? io_r_288_b : _GEN_24067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24069 = 9'h121 == r_count_59_io_out ? io_r_289_b : _GEN_24068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24070 = 9'h122 == r_count_59_io_out ? io_r_290_b : _GEN_24069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24071 = 9'h123 == r_count_59_io_out ? io_r_291_b : _GEN_24070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24072 = 9'h124 == r_count_59_io_out ? io_r_292_b : _GEN_24071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24073 = 9'h125 == r_count_59_io_out ? io_r_293_b : _GEN_24072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24074 = 9'h126 == r_count_59_io_out ? io_r_294_b : _GEN_24073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24075 = 9'h127 == r_count_59_io_out ? io_r_295_b : _GEN_24074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24076 = 9'h128 == r_count_59_io_out ? io_r_296_b : _GEN_24075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24077 = 9'h129 == r_count_59_io_out ? io_r_297_b : _GEN_24076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24078 = 9'h12a == r_count_59_io_out ? io_r_298_b : _GEN_24077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24079 = 9'h12b == r_count_59_io_out ? io_r_299_b : _GEN_24078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24080 = 9'h12c == r_count_59_io_out ? io_r_300_b : _GEN_24079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24081 = 9'h12d == r_count_59_io_out ? io_r_301_b : _GEN_24080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24082 = 9'h12e == r_count_59_io_out ? io_r_302_b : _GEN_24081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24083 = 9'h12f == r_count_59_io_out ? io_r_303_b : _GEN_24082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24084 = 9'h130 == r_count_59_io_out ? io_r_304_b : _GEN_24083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24085 = 9'h131 == r_count_59_io_out ? io_r_305_b : _GEN_24084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24086 = 9'h132 == r_count_59_io_out ? io_r_306_b : _GEN_24085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24087 = 9'h133 == r_count_59_io_out ? io_r_307_b : _GEN_24086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24088 = 9'h134 == r_count_59_io_out ? io_r_308_b : _GEN_24087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24089 = 9'h135 == r_count_59_io_out ? io_r_309_b : _GEN_24088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24090 = 9'h136 == r_count_59_io_out ? io_r_310_b : _GEN_24089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24091 = 9'h137 == r_count_59_io_out ? io_r_311_b : _GEN_24090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24092 = 9'h138 == r_count_59_io_out ? io_r_312_b : _GEN_24091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24093 = 9'h139 == r_count_59_io_out ? io_r_313_b : _GEN_24092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24094 = 9'h13a == r_count_59_io_out ? io_r_314_b : _GEN_24093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24095 = 9'h13b == r_count_59_io_out ? io_r_315_b : _GEN_24094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24096 = 9'h13c == r_count_59_io_out ? io_r_316_b : _GEN_24095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24097 = 9'h13d == r_count_59_io_out ? io_r_317_b : _GEN_24096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24098 = 9'h13e == r_count_59_io_out ? io_r_318_b : _GEN_24097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24099 = 9'h13f == r_count_59_io_out ? io_r_319_b : _GEN_24098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24100 = 9'h140 == r_count_59_io_out ? io_r_320_b : _GEN_24099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24101 = 9'h141 == r_count_59_io_out ? io_r_321_b : _GEN_24100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24102 = 9'h142 == r_count_59_io_out ? io_r_322_b : _GEN_24101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24103 = 9'h143 == r_count_59_io_out ? io_r_323_b : _GEN_24102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24104 = 9'h144 == r_count_59_io_out ? io_r_324_b : _GEN_24103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24105 = 9'h145 == r_count_59_io_out ? io_r_325_b : _GEN_24104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24106 = 9'h146 == r_count_59_io_out ? io_r_326_b : _GEN_24105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24107 = 9'h147 == r_count_59_io_out ? io_r_327_b : _GEN_24106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24108 = 9'h148 == r_count_59_io_out ? io_r_328_b : _GEN_24107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24109 = 9'h149 == r_count_59_io_out ? io_r_329_b : _GEN_24108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24110 = 9'h14a == r_count_59_io_out ? io_r_330_b : _GEN_24109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24111 = 9'h14b == r_count_59_io_out ? io_r_331_b : _GEN_24110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24112 = 9'h14c == r_count_59_io_out ? io_r_332_b : _GEN_24111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24113 = 9'h14d == r_count_59_io_out ? io_r_333_b : _GEN_24112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24114 = 9'h14e == r_count_59_io_out ? io_r_334_b : _GEN_24113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24115 = 9'h14f == r_count_59_io_out ? io_r_335_b : _GEN_24114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24116 = 9'h150 == r_count_59_io_out ? io_r_336_b : _GEN_24115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24117 = 9'h151 == r_count_59_io_out ? io_r_337_b : _GEN_24116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24118 = 9'h152 == r_count_59_io_out ? io_r_338_b : _GEN_24117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24119 = 9'h153 == r_count_59_io_out ? io_r_339_b : _GEN_24118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24120 = 9'h154 == r_count_59_io_out ? io_r_340_b : _GEN_24119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24121 = 9'h155 == r_count_59_io_out ? io_r_341_b : _GEN_24120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24122 = 9'h156 == r_count_59_io_out ? io_r_342_b : _GEN_24121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24123 = 9'h157 == r_count_59_io_out ? io_r_343_b : _GEN_24122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24124 = 9'h158 == r_count_59_io_out ? io_r_344_b : _GEN_24123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24125 = 9'h159 == r_count_59_io_out ? io_r_345_b : _GEN_24124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24126 = 9'h15a == r_count_59_io_out ? io_r_346_b : _GEN_24125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24127 = 9'h15b == r_count_59_io_out ? io_r_347_b : _GEN_24126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24128 = 9'h15c == r_count_59_io_out ? io_r_348_b : _GEN_24127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24129 = 9'h15d == r_count_59_io_out ? io_r_349_b : _GEN_24128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24130 = 9'h15e == r_count_59_io_out ? io_r_350_b : _GEN_24129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24131 = 9'h15f == r_count_59_io_out ? io_r_351_b : _GEN_24130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24132 = 9'h160 == r_count_59_io_out ? io_r_352_b : _GEN_24131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24133 = 9'h161 == r_count_59_io_out ? io_r_353_b : _GEN_24132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24134 = 9'h162 == r_count_59_io_out ? io_r_354_b : _GEN_24133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24135 = 9'h163 == r_count_59_io_out ? io_r_355_b : _GEN_24134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24136 = 9'h164 == r_count_59_io_out ? io_r_356_b : _GEN_24135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24137 = 9'h165 == r_count_59_io_out ? io_r_357_b : _GEN_24136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24138 = 9'h166 == r_count_59_io_out ? io_r_358_b : _GEN_24137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24139 = 9'h167 == r_count_59_io_out ? io_r_359_b : _GEN_24138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24140 = 9'h168 == r_count_59_io_out ? io_r_360_b : _GEN_24139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24141 = 9'h169 == r_count_59_io_out ? io_r_361_b : _GEN_24140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24142 = 9'h16a == r_count_59_io_out ? io_r_362_b : _GEN_24141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24143 = 9'h16b == r_count_59_io_out ? io_r_363_b : _GEN_24142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24144 = 9'h16c == r_count_59_io_out ? io_r_364_b : _GEN_24143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24145 = 9'h16d == r_count_59_io_out ? io_r_365_b : _GEN_24144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24146 = 9'h16e == r_count_59_io_out ? io_r_366_b : _GEN_24145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24147 = 9'h16f == r_count_59_io_out ? io_r_367_b : _GEN_24146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24148 = 9'h170 == r_count_59_io_out ? io_r_368_b : _GEN_24147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24149 = 9'h171 == r_count_59_io_out ? io_r_369_b : _GEN_24148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24150 = 9'h172 == r_count_59_io_out ? io_r_370_b : _GEN_24149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24151 = 9'h173 == r_count_59_io_out ? io_r_371_b : _GEN_24150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24152 = 9'h174 == r_count_59_io_out ? io_r_372_b : _GEN_24151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24153 = 9'h175 == r_count_59_io_out ? io_r_373_b : _GEN_24152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24154 = 9'h176 == r_count_59_io_out ? io_r_374_b : _GEN_24153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24155 = 9'h177 == r_count_59_io_out ? io_r_375_b : _GEN_24154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24156 = 9'h178 == r_count_59_io_out ? io_r_376_b : _GEN_24155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24157 = 9'h179 == r_count_59_io_out ? io_r_377_b : _GEN_24156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24158 = 9'h17a == r_count_59_io_out ? io_r_378_b : _GEN_24157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24159 = 9'h17b == r_count_59_io_out ? io_r_379_b : _GEN_24158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24160 = 9'h17c == r_count_59_io_out ? io_r_380_b : _GEN_24159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24161 = 9'h17d == r_count_59_io_out ? io_r_381_b : _GEN_24160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24162 = 9'h17e == r_count_59_io_out ? io_r_382_b : _GEN_24161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24163 = 9'h17f == r_count_59_io_out ? io_r_383_b : _GEN_24162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24164 = 9'h180 == r_count_59_io_out ? io_r_384_b : _GEN_24163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24165 = 9'h181 == r_count_59_io_out ? io_r_385_b : _GEN_24164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24166 = 9'h182 == r_count_59_io_out ? io_r_386_b : _GEN_24165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24167 = 9'h183 == r_count_59_io_out ? io_r_387_b : _GEN_24166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24168 = 9'h184 == r_count_59_io_out ? io_r_388_b : _GEN_24167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24169 = 9'h185 == r_count_59_io_out ? io_r_389_b : _GEN_24168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24170 = 9'h186 == r_count_59_io_out ? io_r_390_b : _GEN_24169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24171 = 9'h187 == r_count_59_io_out ? io_r_391_b : _GEN_24170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24172 = 9'h188 == r_count_59_io_out ? io_r_392_b : _GEN_24171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24173 = 9'h189 == r_count_59_io_out ? io_r_393_b : _GEN_24172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24174 = 9'h18a == r_count_59_io_out ? io_r_394_b : _GEN_24173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24175 = 9'h18b == r_count_59_io_out ? io_r_395_b : _GEN_24174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24176 = 9'h18c == r_count_59_io_out ? io_r_396_b : _GEN_24175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24177 = 9'h18d == r_count_59_io_out ? io_r_397_b : _GEN_24176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_24178 = 9'h18e == r_count_59_io_out ? io_r_398_b : _GEN_24177; // @[SWChisel.scala 221:{19,19}]
  SWCell array_0 ( // @[SWChisel.scala 170:39]
    .io_q(array_0_io_q),
    .io_r(array_0_io_r),
    .io_e_i(array_0_io_e_i),
    .io_f_i(array_0_io_f_i),
    .io_ve_i(array_0_io_ve_i),
    .io_vf_i(array_0_io_vf_i),
    .io_vv_i(array_0_io_vv_i),
    .io_e_o(array_0_io_e_o),
    .io_f_o(array_0_io_f_o),
    .io_v_o(array_0_io_v_o)
  );
  SWCell array_1 ( // @[SWChisel.scala 170:39]
    .io_q(array_1_io_q),
    .io_r(array_1_io_r),
    .io_e_i(array_1_io_e_i),
    .io_f_i(array_1_io_f_i),
    .io_ve_i(array_1_io_ve_i),
    .io_vf_i(array_1_io_vf_i),
    .io_vv_i(array_1_io_vv_i),
    .io_e_o(array_1_io_e_o),
    .io_f_o(array_1_io_f_o),
    .io_v_o(array_1_io_v_o)
  );
  SWCell array_2 ( // @[SWChisel.scala 170:39]
    .io_q(array_2_io_q),
    .io_r(array_2_io_r),
    .io_e_i(array_2_io_e_i),
    .io_f_i(array_2_io_f_i),
    .io_ve_i(array_2_io_ve_i),
    .io_vf_i(array_2_io_vf_i),
    .io_vv_i(array_2_io_vv_i),
    .io_e_o(array_2_io_e_o),
    .io_f_o(array_2_io_f_o),
    .io_v_o(array_2_io_v_o)
  );
  SWCell array_3 ( // @[SWChisel.scala 170:39]
    .io_q(array_3_io_q),
    .io_r(array_3_io_r),
    .io_e_i(array_3_io_e_i),
    .io_f_i(array_3_io_f_i),
    .io_ve_i(array_3_io_ve_i),
    .io_vf_i(array_3_io_vf_i),
    .io_vv_i(array_3_io_vv_i),
    .io_e_o(array_3_io_e_o),
    .io_f_o(array_3_io_f_o),
    .io_v_o(array_3_io_v_o)
  );
  SWCell array_4 ( // @[SWChisel.scala 170:39]
    .io_q(array_4_io_q),
    .io_r(array_4_io_r),
    .io_e_i(array_4_io_e_i),
    .io_f_i(array_4_io_f_i),
    .io_ve_i(array_4_io_ve_i),
    .io_vf_i(array_4_io_vf_i),
    .io_vv_i(array_4_io_vv_i),
    .io_e_o(array_4_io_e_o),
    .io_f_o(array_4_io_f_o),
    .io_v_o(array_4_io_v_o)
  );
  SWCell array_5 ( // @[SWChisel.scala 170:39]
    .io_q(array_5_io_q),
    .io_r(array_5_io_r),
    .io_e_i(array_5_io_e_i),
    .io_f_i(array_5_io_f_i),
    .io_ve_i(array_5_io_ve_i),
    .io_vf_i(array_5_io_vf_i),
    .io_vv_i(array_5_io_vv_i),
    .io_e_o(array_5_io_e_o),
    .io_f_o(array_5_io_f_o),
    .io_v_o(array_5_io_v_o)
  );
  SWCell array_6 ( // @[SWChisel.scala 170:39]
    .io_q(array_6_io_q),
    .io_r(array_6_io_r),
    .io_e_i(array_6_io_e_i),
    .io_f_i(array_6_io_f_i),
    .io_ve_i(array_6_io_ve_i),
    .io_vf_i(array_6_io_vf_i),
    .io_vv_i(array_6_io_vv_i),
    .io_e_o(array_6_io_e_o),
    .io_f_o(array_6_io_f_o),
    .io_v_o(array_6_io_v_o)
  );
  SWCell array_7 ( // @[SWChisel.scala 170:39]
    .io_q(array_7_io_q),
    .io_r(array_7_io_r),
    .io_e_i(array_7_io_e_i),
    .io_f_i(array_7_io_f_i),
    .io_ve_i(array_7_io_ve_i),
    .io_vf_i(array_7_io_vf_i),
    .io_vv_i(array_7_io_vv_i),
    .io_e_o(array_7_io_e_o),
    .io_f_o(array_7_io_f_o),
    .io_v_o(array_7_io_v_o)
  );
  SWCell array_8 ( // @[SWChisel.scala 170:39]
    .io_q(array_8_io_q),
    .io_r(array_8_io_r),
    .io_e_i(array_8_io_e_i),
    .io_f_i(array_8_io_f_i),
    .io_ve_i(array_8_io_ve_i),
    .io_vf_i(array_8_io_vf_i),
    .io_vv_i(array_8_io_vv_i),
    .io_e_o(array_8_io_e_o),
    .io_f_o(array_8_io_f_o),
    .io_v_o(array_8_io_v_o)
  );
  SWCell array_9 ( // @[SWChisel.scala 170:39]
    .io_q(array_9_io_q),
    .io_r(array_9_io_r),
    .io_e_i(array_9_io_e_i),
    .io_f_i(array_9_io_f_i),
    .io_ve_i(array_9_io_ve_i),
    .io_vf_i(array_9_io_vf_i),
    .io_vv_i(array_9_io_vv_i),
    .io_e_o(array_9_io_e_o),
    .io_f_o(array_9_io_f_o),
    .io_v_o(array_9_io_v_o)
  );
  SWCell array_10 ( // @[SWChisel.scala 170:39]
    .io_q(array_10_io_q),
    .io_r(array_10_io_r),
    .io_e_i(array_10_io_e_i),
    .io_f_i(array_10_io_f_i),
    .io_ve_i(array_10_io_ve_i),
    .io_vf_i(array_10_io_vf_i),
    .io_vv_i(array_10_io_vv_i),
    .io_e_o(array_10_io_e_o),
    .io_f_o(array_10_io_f_o),
    .io_v_o(array_10_io_v_o)
  );
  SWCell array_11 ( // @[SWChisel.scala 170:39]
    .io_q(array_11_io_q),
    .io_r(array_11_io_r),
    .io_e_i(array_11_io_e_i),
    .io_f_i(array_11_io_f_i),
    .io_ve_i(array_11_io_ve_i),
    .io_vf_i(array_11_io_vf_i),
    .io_vv_i(array_11_io_vv_i),
    .io_e_o(array_11_io_e_o),
    .io_f_o(array_11_io_f_o),
    .io_v_o(array_11_io_v_o)
  );
  SWCell array_12 ( // @[SWChisel.scala 170:39]
    .io_q(array_12_io_q),
    .io_r(array_12_io_r),
    .io_e_i(array_12_io_e_i),
    .io_f_i(array_12_io_f_i),
    .io_ve_i(array_12_io_ve_i),
    .io_vf_i(array_12_io_vf_i),
    .io_vv_i(array_12_io_vv_i),
    .io_e_o(array_12_io_e_o),
    .io_f_o(array_12_io_f_o),
    .io_v_o(array_12_io_v_o)
  );
  SWCell array_13 ( // @[SWChisel.scala 170:39]
    .io_q(array_13_io_q),
    .io_r(array_13_io_r),
    .io_e_i(array_13_io_e_i),
    .io_f_i(array_13_io_f_i),
    .io_ve_i(array_13_io_ve_i),
    .io_vf_i(array_13_io_vf_i),
    .io_vv_i(array_13_io_vv_i),
    .io_e_o(array_13_io_e_o),
    .io_f_o(array_13_io_f_o),
    .io_v_o(array_13_io_v_o)
  );
  SWCell array_14 ( // @[SWChisel.scala 170:39]
    .io_q(array_14_io_q),
    .io_r(array_14_io_r),
    .io_e_i(array_14_io_e_i),
    .io_f_i(array_14_io_f_i),
    .io_ve_i(array_14_io_ve_i),
    .io_vf_i(array_14_io_vf_i),
    .io_vv_i(array_14_io_vv_i),
    .io_e_o(array_14_io_e_o),
    .io_f_o(array_14_io_f_o),
    .io_v_o(array_14_io_v_o)
  );
  SWCell array_15 ( // @[SWChisel.scala 170:39]
    .io_q(array_15_io_q),
    .io_r(array_15_io_r),
    .io_e_i(array_15_io_e_i),
    .io_f_i(array_15_io_f_i),
    .io_ve_i(array_15_io_ve_i),
    .io_vf_i(array_15_io_vf_i),
    .io_vv_i(array_15_io_vv_i),
    .io_e_o(array_15_io_e_o),
    .io_f_o(array_15_io_f_o),
    .io_v_o(array_15_io_v_o)
  );
  SWCell array_16 ( // @[SWChisel.scala 170:39]
    .io_q(array_16_io_q),
    .io_r(array_16_io_r),
    .io_e_i(array_16_io_e_i),
    .io_f_i(array_16_io_f_i),
    .io_ve_i(array_16_io_ve_i),
    .io_vf_i(array_16_io_vf_i),
    .io_vv_i(array_16_io_vv_i),
    .io_e_o(array_16_io_e_o),
    .io_f_o(array_16_io_f_o),
    .io_v_o(array_16_io_v_o)
  );
  SWCell array_17 ( // @[SWChisel.scala 170:39]
    .io_q(array_17_io_q),
    .io_r(array_17_io_r),
    .io_e_i(array_17_io_e_i),
    .io_f_i(array_17_io_f_i),
    .io_ve_i(array_17_io_ve_i),
    .io_vf_i(array_17_io_vf_i),
    .io_vv_i(array_17_io_vv_i),
    .io_e_o(array_17_io_e_o),
    .io_f_o(array_17_io_f_o),
    .io_v_o(array_17_io_v_o)
  );
  SWCell array_18 ( // @[SWChisel.scala 170:39]
    .io_q(array_18_io_q),
    .io_r(array_18_io_r),
    .io_e_i(array_18_io_e_i),
    .io_f_i(array_18_io_f_i),
    .io_ve_i(array_18_io_ve_i),
    .io_vf_i(array_18_io_vf_i),
    .io_vv_i(array_18_io_vv_i),
    .io_e_o(array_18_io_e_o),
    .io_f_o(array_18_io_f_o),
    .io_v_o(array_18_io_v_o)
  );
  SWCell array_19 ( // @[SWChisel.scala 170:39]
    .io_q(array_19_io_q),
    .io_r(array_19_io_r),
    .io_e_i(array_19_io_e_i),
    .io_f_i(array_19_io_f_i),
    .io_ve_i(array_19_io_ve_i),
    .io_vf_i(array_19_io_vf_i),
    .io_vv_i(array_19_io_vv_i),
    .io_e_o(array_19_io_e_o),
    .io_f_o(array_19_io_f_o),
    .io_v_o(array_19_io_v_o)
  );
  SWCell array_20 ( // @[SWChisel.scala 170:39]
    .io_q(array_20_io_q),
    .io_r(array_20_io_r),
    .io_e_i(array_20_io_e_i),
    .io_f_i(array_20_io_f_i),
    .io_ve_i(array_20_io_ve_i),
    .io_vf_i(array_20_io_vf_i),
    .io_vv_i(array_20_io_vv_i),
    .io_e_o(array_20_io_e_o),
    .io_f_o(array_20_io_f_o),
    .io_v_o(array_20_io_v_o)
  );
  SWCell array_21 ( // @[SWChisel.scala 170:39]
    .io_q(array_21_io_q),
    .io_r(array_21_io_r),
    .io_e_i(array_21_io_e_i),
    .io_f_i(array_21_io_f_i),
    .io_ve_i(array_21_io_ve_i),
    .io_vf_i(array_21_io_vf_i),
    .io_vv_i(array_21_io_vv_i),
    .io_e_o(array_21_io_e_o),
    .io_f_o(array_21_io_f_o),
    .io_v_o(array_21_io_v_o)
  );
  SWCell array_22 ( // @[SWChisel.scala 170:39]
    .io_q(array_22_io_q),
    .io_r(array_22_io_r),
    .io_e_i(array_22_io_e_i),
    .io_f_i(array_22_io_f_i),
    .io_ve_i(array_22_io_ve_i),
    .io_vf_i(array_22_io_vf_i),
    .io_vv_i(array_22_io_vv_i),
    .io_e_o(array_22_io_e_o),
    .io_f_o(array_22_io_f_o),
    .io_v_o(array_22_io_v_o)
  );
  SWCell array_23 ( // @[SWChisel.scala 170:39]
    .io_q(array_23_io_q),
    .io_r(array_23_io_r),
    .io_e_i(array_23_io_e_i),
    .io_f_i(array_23_io_f_i),
    .io_ve_i(array_23_io_ve_i),
    .io_vf_i(array_23_io_vf_i),
    .io_vv_i(array_23_io_vv_i),
    .io_e_o(array_23_io_e_o),
    .io_f_o(array_23_io_f_o),
    .io_v_o(array_23_io_v_o)
  );
  SWCell array_24 ( // @[SWChisel.scala 170:39]
    .io_q(array_24_io_q),
    .io_r(array_24_io_r),
    .io_e_i(array_24_io_e_i),
    .io_f_i(array_24_io_f_i),
    .io_ve_i(array_24_io_ve_i),
    .io_vf_i(array_24_io_vf_i),
    .io_vv_i(array_24_io_vv_i),
    .io_e_o(array_24_io_e_o),
    .io_f_o(array_24_io_f_o),
    .io_v_o(array_24_io_v_o)
  );
  SWCell array_25 ( // @[SWChisel.scala 170:39]
    .io_q(array_25_io_q),
    .io_r(array_25_io_r),
    .io_e_i(array_25_io_e_i),
    .io_f_i(array_25_io_f_i),
    .io_ve_i(array_25_io_ve_i),
    .io_vf_i(array_25_io_vf_i),
    .io_vv_i(array_25_io_vv_i),
    .io_e_o(array_25_io_e_o),
    .io_f_o(array_25_io_f_o),
    .io_v_o(array_25_io_v_o)
  );
  SWCell array_26 ( // @[SWChisel.scala 170:39]
    .io_q(array_26_io_q),
    .io_r(array_26_io_r),
    .io_e_i(array_26_io_e_i),
    .io_f_i(array_26_io_f_i),
    .io_ve_i(array_26_io_ve_i),
    .io_vf_i(array_26_io_vf_i),
    .io_vv_i(array_26_io_vv_i),
    .io_e_o(array_26_io_e_o),
    .io_f_o(array_26_io_f_o),
    .io_v_o(array_26_io_v_o)
  );
  SWCell array_27 ( // @[SWChisel.scala 170:39]
    .io_q(array_27_io_q),
    .io_r(array_27_io_r),
    .io_e_i(array_27_io_e_i),
    .io_f_i(array_27_io_f_i),
    .io_ve_i(array_27_io_ve_i),
    .io_vf_i(array_27_io_vf_i),
    .io_vv_i(array_27_io_vv_i),
    .io_e_o(array_27_io_e_o),
    .io_f_o(array_27_io_f_o),
    .io_v_o(array_27_io_v_o)
  );
  SWCell array_28 ( // @[SWChisel.scala 170:39]
    .io_q(array_28_io_q),
    .io_r(array_28_io_r),
    .io_e_i(array_28_io_e_i),
    .io_f_i(array_28_io_f_i),
    .io_ve_i(array_28_io_ve_i),
    .io_vf_i(array_28_io_vf_i),
    .io_vv_i(array_28_io_vv_i),
    .io_e_o(array_28_io_e_o),
    .io_f_o(array_28_io_f_o),
    .io_v_o(array_28_io_v_o)
  );
  SWCell array_29 ( // @[SWChisel.scala 170:39]
    .io_q(array_29_io_q),
    .io_r(array_29_io_r),
    .io_e_i(array_29_io_e_i),
    .io_f_i(array_29_io_f_i),
    .io_ve_i(array_29_io_ve_i),
    .io_vf_i(array_29_io_vf_i),
    .io_vv_i(array_29_io_vv_i),
    .io_e_o(array_29_io_e_o),
    .io_f_o(array_29_io_f_o),
    .io_v_o(array_29_io_v_o)
  );
  SWCell array_30 ( // @[SWChisel.scala 170:39]
    .io_q(array_30_io_q),
    .io_r(array_30_io_r),
    .io_e_i(array_30_io_e_i),
    .io_f_i(array_30_io_f_i),
    .io_ve_i(array_30_io_ve_i),
    .io_vf_i(array_30_io_vf_i),
    .io_vv_i(array_30_io_vv_i),
    .io_e_o(array_30_io_e_o),
    .io_f_o(array_30_io_f_o),
    .io_v_o(array_30_io_v_o)
  );
  SWCell array_31 ( // @[SWChisel.scala 170:39]
    .io_q(array_31_io_q),
    .io_r(array_31_io_r),
    .io_e_i(array_31_io_e_i),
    .io_f_i(array_31_io_f_i),
    .io_ve_i(array_31_io_ve_i),
    .io_vf_i(array_31_io_vf_i),
    .io_vv_i(array_31_io_vv_i),
    .io_e_o(array_31_io_e_o),
    .io_f_o(array_31_io_f_o),
    .io_v_o(array_31_io_v_o)
  );
  SWCell array_32 ( // @[SWChisel.scala 170:39]
    .io_q(array_32_io_q),
    .io_r(array_32_io_r),
    .io_e_i(array_32_io_e_i),
    .io_f_i(array_32_io_f_i),
    .io_ve_i(array_32_io_ve_i),
    .io_vf_i(array_32_io_vf_i),
    .io_vv_i(array_32_io_vv_i),
    .io_e_o(array_32_io_e_o),
    .io_f_o(array_32_io_f_o),
    .io_v_o(array_32_io_v_o)
  );
  SWCell array_33 ( // @[SWChisel.scala 170:39]
    .io_q(array_33_io_q),
    .io_r(array_33_io_r),
    .io_e_i(array_33_io_e_i),
    .io_f_i(array_33_io_f_i),
    .io_ve_i(array_33_io_ve_i),
    .io_vf_i(array_33_io_vf_i),
    .io_vv_i(array_33_io_vv_i),
    .io_e_o(array_33_io_e_o),
    .io_f_o(array_33_io_f_o),
    .io_v_o(array_33_io_v_o)
  );
  SWCell array_34 ( // @[SWChisel.scala 170:39]
    .io_q(array_34_io_q),
    .io_r(array_34_io_r),
    .io_e_i(array_34_io_e_i),
    .io_f_i(array_34_io_f_i),
    .io_ve_i(array_34_io_ve_i),
    .io_vf_i(array_34_io_vf_i),
    .io_vv_i(array_34_io_vv_i),
    .io_e_o(array_34_io_e_o),
    .io_f_o(array_34_io_f_o),
    .io_v_o(array_34_io_v_o)
  );
  SWCell array_35 ( // @[SWChisel.scala 170:39]
    .io_q(array_35_io_q),
    .io_r(array_35_io_r),
    .io_e_i(array_35_io_e_i),
    .io_f_i(array_35_io_f_i),
    .io_ve_i(array_35_io_ve_i),
    .io_vf_i(array_35_io_vf_i),
    .io_vv_i(array_35_io_vv_i),
    .io_e_o(array_35_io_e_o),
    .io_f_o(array_35_io_f_o),
    .io_v_o(array_35_io_v_o)
  );
  SWCell array_36 ( // @[SWChisel.scala 170:39]
    .io_q(array_36_io_q),
    .io_r(array_36_io_r),
    .io_e_i(array_36_io_e_i),
    .io_f_i(array_36_io_f_i),
    .io_ve_i(array_36_io_ve_i),
    .io_vf_i(array_36_io_vf_i),
    .io_vv_i(array_36_io_vv_i),
    .io_e_o(array_36_io_e_o),
    .io_f_o(array_36_io_f_o),
    .io_v_o(array_36_io_v_o)
  );
  SWCell array_37 ( // @[SWChisel.scala 170:39]
    .io_q(array_37_io_q),
    .io_r(array_37_io_r),
    .io_e_i(array_37_io_e_i),
    .io_f_i(array_37_io_f_i),
    .io_ve_i(array_37_io_ve_i),
    .io_vf_i(array_37_io_vf_i),
    .io_vv_i(array_37_io_vv_i),
    .io_e_o(array_37_io_e_o),
    .io_f_o(array_37_io_f_o),
    .io_v_o(array_37_io_v_o)
  );
  SWCell array_38 ( // @[SWChisel.scala 170:39]
    .io_q(array_38_io_q),
    .io_r(array_38_io_r),
    .io_e_i(array_38_io_e_i),
    .io_f_i(array_38_io_f_i),
    .io_ve_i(array_38_io_ve_i),
    .io_vf_i(array_38_io_vf_i),
    .io_vv_i(array_38_io_vv_i),
    .io_e_o(array_38_io_e_o),
    .io_f_o(array_38_io_f_o),
    .io_v_o(array_38_io_v_o)
  );
  SWCell array_39 ( // @[SWChisel.scala 170:39]
    .io_q(array_39_io_q),
    .io_r(array_39_io_r),
    .io_e_i(array_39_io_e_i),
    .io_f_i(array_39_io_f_i),
    .io_ve_i(array_39_io_ve_i),
    .io_vf_i(array_39_io_vf_i),
    .io_vv_i(array_39_io_vv_i),
    .io_e_o(array_39_io_e_o),
    .io_f_o(array_39_io_f_o),
    .io_v_o(array_39_io_v_o)
  );
  SWCell array_40 ( // @[SWChisel.scala 170:39]
    .io_q(array_40_io_q),
    .io_r(array_40_io_r),
    .io_e_i(array_40_io_e_i),
    .io_f_i(array_40_io_f_i),
    .io_ve_i(array_40_io_ve_i),
    .io_vf_i(array_40_io_vf_i),
    .io_vv_i(array_40_io_vv_i),
    .io_e_o(array_40_io_e_o),
    .io_f_o(array_40_io_f_o),
    .io_v_o(array_40_io_v_o)
  );
  SWCell array_41 ( // @[SWChisel.scala 170:39]
    .io_q(array_41_io_q),
    .io_r(array_41_io_r),
    .io_e_i(array_41_io_e_i),
    .io_f_i(array_41_io_f_i),
    .io_ve_i(array_41_io_ve_i),
    .io_vf_i(array_41_io_vf_i),
    .io_vv_i(array_41_io_vv_i),
    .io_e_o(array_41_io_e_o),
    .io_f_o(array_41_io_f_o),
    .io_v_o(array_41_io_v_o)
  );
  SWCell array_42 ( // @[SWChisel.scala 170:39]
    .io_q(array_42_io_q),
    .io_r(array_42_io_r),
    .io_e_i(array_42_io_e_i),
    .io_f_i(array_42_io_f_i),
    .io_ve_i(array_42_io_ve_i),
    .io_vf_i(array_42_io_vf_i),
    .io_vv_i(array_42_io_vv_i),
    .io_e_o(array_42_io_e_o),
    .io_f_o(array_42_io_f_o),
    .io_v_o(array_42_io_v_o)
  );
  SWCell array_43 ( // @[SWChisel.scala 170:39]
    .io_q(array_43_io_q),
    .io_r(array_43_io_r),
    .io_e_i(array_43_io_e_i),
    .io_f_i(array_43_io_f_i),
    .io_ve_i(array_43_io_ve_i),
    .io_vf_i(array_43_io_vf_i),
    .io_vv_i(array_43_io_vv_i),
    .io_e_o(array_43_io_e_o),
    .io_f_o(array_43_io_f_o),
    .io_v_o(array_43_io_v_o)
  );
  SWCell array_44 ( // @[SWChisel.scala 170:39]
    .io_q(array_44_io_q),
    .io_r(array_44_io_r),
    .io_e_i(array_44_io_e_i),
    .io_f_i(array_44_io_f_i),
    .io_ve_i(array_44_io_ve_i),
    .io_vf_i(array_44_io_vf_i),
    .io_vv_i(array_44_io_vv_i),
    .io_e_o(array_44_io_e_o),
    .io_f_o(array_44_io_f_o),
    .io_v_o(array_44_io_v_o)
  );
  SWCell array_45 ( // @[SWChisel.scala 170:39]
    .io_q(array_45_io_q),
    .io_r(array_45_io_r),
    .io_e_i(array_45_io_e_i),
    .io_f_i(array_45_io_f_i),
    .io_ve_i(array_45_io_ve_i),
    .io_vf_i(array_45_io_vf_i),
    .io_vv_i(array_45_io_vv_i),
    .io_e_o(array_45_io_e_o),
    .io_f_o(array_45_io_f_o),
    .io_v_o(array_45_io_v_o)
  );
  SWCell array_46 ( // @[SWChisel.scala 170:39]
    .io_q(array_46_io_q),
    .io_r(array_46_io_r),
    .io_e_i(array_46_io_e_i),
    .io_f_i(array_46_io_f_i),
    .io_ve_i(array_46_io_ve_i),
    .io_vf_i(array_46_io_vf_i),
    .io_vv_i(array_46_io_vv_i),
    .io_e_o(array_46_io_e_o),
    .io_f_o(array_46_io_f_o),
    .io_v_o(array_46_io_v_o)
  );
  SWCell array_47 ( // @[SWChisel.scala 170:39]
    .io_q(array_47_io_q),
    .io_r(array_47_io_r),
    .io_e_i(array_47_io_e_i),
    .io_f_i(array_47_io_f_i),
    .io_ve_i(array_47_io_ve_i),
    .io_vf_i(array_47_io_vf_i),
    .io_vv_i(array_47_io_vv_i),
    .io_e_o(array_47_io_e_o),
    .io_f_o(array_47_io_f_o),
    .io_v_o(array_47_io_v_o)
  );
  SWCell array_48 ( // @[SWChisel.scala 170:39]
    .io_q(array_48_io_q),
    .io_r(array_48_io_r),
    .io_e_i(array_48_io_e_i),
    .io_f_i(array_48_io_f_i),
    .io_ve_i(array_48_io_ve_i),
    .io_vf_i(array_48_io_vf_i),
    .io_vv_i(array_48_io_vv_i),
    .io_e_o(array_48_io_e_o),
    .io_f_o(array_48_io_f_o),
    .io_v_o(array_48_io_v_o)
  );
  SWCell array_49 ( // @[SWChisel.scala 170:39]
    .io_q(array_49_io_q),
    .io_r(array_49_io_r),
    .io_e_i(array_49_io_e_i),
    .io_f_i(array_49_io_f_i),
    .io_ve_i(array_49_io_ve_i),
    .io_vf_i(array_49_io_vf_i),
    .io_vv_i(array_49_io_vv_i),
    .io_e_o(array_49_io_e_o),
    .io_f_o(array_49_io_f_o),
    .io_v_o(array_49_io_v_o)
  );
  SWCell array_50 ( // @[SWChisel.scala 170:39]
    .io_q(array_50_io_q),
    .io_r(array_50_io_r),
    .io_e_i(array_50_io_e_i),
    .io_f_i(array_50_io_f_i),
    .io_ve_i(array_50_io_ve_i),
    .io_vf_i(array_50_io_vf_i),
    .io_vv_i(array_50_io_vv_i),
    .io_e_o(array_50_io_e_o),
    .io_f_o(array_50_io_f_o),
    .io_v_o(array_50_io_v_o)
  );
  SWCell array_51 ( // @[SWChisel.scala 170:39]
    .io_q(array_51_io_q),
    .io_r(array_51_io_r),
    .io_e_i(array_51_io_e_i),
    .io_f_i(array_51_io_f_i),
    .io_ve_i(array_51_io_ve_i),
    .io_vf_i(array_51_io_vf_i),
    .io_vv_i(array_51_io_vv_i),
    .io_e_o(array_51_io_e_o),
    .io_f_o(array_51_io_f_o),
    .io_v_o(array_51_io_v_o)
  );
  SWCell array_52 ( // @[SWChisel.scala 170:39]
    .io_q(array_52_io_q),
    .io_r(array_52_io_r),
    .io_e_i(array_52_io_e_i),
    .io_f_i(array_52_io_f_i),
    .io_ve_i(array_52_io_ve_i),
    .io_vf_i(array_52_io_vf_i),
    .io_vv_i(array_52_io_vv_i),
    .io_e_o(array_52_io_e_o),
    .io_f_o(array_52_io_f_o),
    .io_v_o(array_52_io_v_o)
  );
  SWCell array_53 ( // @[SWChisel.scala 170:39]
    .io_q(array_53_io_q),
    .io_r(array_53_io_r),
    .io_e_i(array_53_io_e_i),
    .io_f_i(array_53_io_f_i),
    .io_ve_i(array_53_io_ve_i),
    .io_vf_i(array_53_io_vf_i),
    .io_vv_i(array_53_io_vv_i),
    .io_e_o(array_53_io_e_o),
    .io_f_o(array_53_io_f_o),
    .io_v_o(array_53_io_v_o)
  );
  SWCell array_54 ( // @[SWChisel.scala 170:39]
    .io_q(array_54_io_q),
    .io_r(array_54_io_r),
    .io_e_i(array_54_io_e_i),
    .io_f_i(array_54_io_f_i),
    .io_ve_i(array_54_io_ve_i),
    .io_vf_i(array_54_io_vf_i),
    .io_vv_i(array_54_io_vv_i),
    .io_e_o(array_54_io_e_o),
    .io_f_o(array_54_io_f_o),
    .io_v_o(array_54_io_v_o)
  );
  SWCell array_55 ( // @[SWChisel.scala 170:39]
    .io_q(array_55_io_q),
    .io_r(array_55_io_r),
    .io_e_i(array_55_io_e_i),
    .io_f_i(array_55_io_f_i),
    .io_ve_i(array_55_io_ve_i),
    .io_vf_i(array_55_io_vf_i),
    .io_vv_i(array_55_io_vv_i),
    .io_e_o(array_55_io_e_o),
    .io_f_o(array_55_io_f_o),
    .io_v_o(array_55_io_v_o)
  );
  SWCell array_56 ( // @[SWChisel.scala 170:39]
    .io_q(array_56_io_q),
    .io_r(array_56_io_r),
    .io_e_i(array_56_io_e_i),
    .io_f_i(array_56_io_f_i),
    .io_ve_i(array_56_io_ve_i),
    .io_vf_i(array_56_io_vf_i),
    .io_vv_i(array_56_io_vv_i),
    .io_e_o(array_56_io_e_o),
    .io_f_o(array_56_io_f_o),
    .io_v_o(array_56_io_v_o)
  );
  SWCell array_57 ( // @[SWChisel.scala 170:39]
    .io_q(array_57_io_q),
    .io_r(array_57_io_r),
    .io_e_i(array_57_io_e_i),
    .io_f_i(array_57_io_f_i),
    .io_ve_i(array_57_io_ve_i),
    .io_vf_i(array_57_io_vf_i),
    .io_vv_i(array_57_io_vv_i),
    .io_e_o(array_57_io_e_o),
    .io_f_o(array_57_io_f_o),
    .io_v_o(array_57_io_v_o)
  );
  SWCell array_58 ( // @[SWChisel.scala 170:39]
    .io_q(array_58_io_q),
    .io_r(array_58_io_r),
    .io_e_i(array_58_io_e_i),
    .io_f_i(array_58_io_f_i),
    .io_ve_i(array_58_io_ve_i),
    .io_vf_i(array_58_io_vf_i),
    .io_vv_i(array_58_io_vv_i),
    .io_e_o(array_58_io_e_o),
    .io_f_o(array_58_io_f_o),
    .io_v_o(array_58_io_v_o)
  );
  SWCell array_59 ( // @[SWChisel.scala 170:39]
    .io_q(array_59_io_q),
    .io_r(array_59_io_r),
    .io_e_i(array_59_io_e_i),
    .io_f_i(array_59_io_f_i),
    .io_ve_i(array_59_io_ve_i),
    .io_vf_i(array_59_io_vf_i),
    .io_vv_i(array_59_io_vv_i),
    .io_e_o(array_59_io_e_o),
    .io_f_o(array_59_io_f_o),
    .io_v_o(array_59_io_v_o)
  );
  MyCounter r_count_0 ( // @[SWChisel.scala 171:41]
    .clock(r_count_0_clock),
    .reset(r_count_0_reset),
    .io_en(r_count_0_io_en),
    .io_out(r_count_0_io_out)
  );
  MyCounter r_count_1 ( // @[SWChisel.scala 171:41]
    .clock(r_count_1_clock),
    .reset(r_count_1_reset),
    .io_en(r_count_1_io_en),
    .io_out(r_count_1_io_out)
  );
  MyCounter r_count_2 ( // @[SWChisel.scala 171:41]
    .clock(r_count_2_clock),
    .reset(r_count_2_reset),
    .io_en(r_count_2_io_en),
    .io_out(r_count_2_io_out)
  );
  MyCounter r_count_3 ( // @[SWChisel.scala 171:41]
    .clock(r_count_3_clock),
    .reset(r_count_3_reset),
    .io_en(r_count_3_io_en),
    .io_out(r_count_3_io_out)
  );
  MyCounter r_count_4 ( // @[SWChisel.scala 171:41]
    .clock(r_count_4_clock),
    .reset(r_count_4_reset),
    .io_en(r_count_4_io_en),
    .io_out(r_count_4_io_out)
  );
  MyCounter r_count_5 ( // @[SWChisel.scala 171:41]
    .clock(r_count_5_clock),
    .reset(r_count_5_reset),
    .io_en(r_count_5_io_en),
    .io_out(r_count_5_io_out)
  );
  MyCounter r_count_6 ( // @[SWChisel.scala 171:41]
    .clock(r_count_6_clock),
    .reset(r_count_6_reset),
    .io_en(r_count_6_io_en),
    .io_out(r_count_6_io_out)
  );
  MyCounter r_count_7 ( // @[SWChisel.scala 171:41]
    .clock(r_count_7_clock),
    .reset(r_count_7_reset),
    .io_en(r_count_7_io_en),
    .io_out(r_count_7_io_out)
  );
  MyCounter r_count_8 ( // @[SWChisel.scala 171:41]
    .clock(r_count_8_clock),
    .reset(r_count_8_reset),
    .io_en(r_count_8_io_en),
    .io_out(r_count_8_io_out)
  );
  MyCounter r_count_9 ( // @[SWChisel.scala 171:41]
    .clock(r_count_9_clock),
    .reset(r_count_9_reset),
    .io_en(r_count_9_io_en),
    .io_out(r_count_9_io_out)
  );
  MyCounter r_count_10 ( // @[SWChisel.scala 171:41]
    .clock(r_count_10_clock),
    .reset(r_count_10_reset),
    .io_en(r_count_10_io_en),
    .io_out(r_count_10_io_out)
  );
  MyCounter r_count_11 ( // @[SWChisel.scala 171:41]
    .clock(r_count_11_clock),
    .reset(r_count_11_reset),
    .io_en(r_count_11_io_en),
    .io_out(r_count_11_io_out)
  );
  MyCounter r_count_12 ( // @[SWChisel.scala 171:41]
    .clock(r_count_12_clock),
    .reset(r_count_12_reset),
    .io_en(r_count_12_io_en),
    .io_out(r_count_12_io_out)
  );
  MyCounter r_count_13 ( // @[SWChisel.scala 171:41]
    .clock(r_count_13_clock),
    .reset(r_count_13_reset),
    .io_en(r_count_13_io_en),
    .io_out(r_count_13_io_out)
  );
  MyCounter r_count_14 ( // @[SWChisel.scala 171:41]
    .clock(r_count_14_clock),
    .reset(r_count_14_reset),
    .io_en(r_count_14_io_en),
    .io_out(r_count_14_io_out)
  );
  MyCounter r_count_15 ( // @[SWChisel.scala 171:41]
    .clock(r_count_15_clock),
    .reset(r_count_15_reset),
    .io_en(r_count_15_io_en),
    .io_out(r_count_15_io_out)
  );
  MyCounter r_count_16 ( // @[SWChisel.scala 171:41]
    .clock(r_count_16_clock),
    .reset(r_count_16_reset),
    .io_en(r_count_16_io_en),
    .io_out(r_count_16_io_out)
  );
  MyCounter r_count_17 ( // @[SWChisel.scala 171:41]
    .clock(r_count_17_clock),
    .reset(r_count_17_reset),
    .io_en(r_count_17_io_en),
    .io_out(r_count_17_io_out)
  );
  MyCounter r_count_18 ( // @[SWChisel.scala 171:41]
    .clock(r_count_18_clock),
    .reset(r_count_18_reset),
    .io_en(r_count_18_io_en),
    .io_out(r_count_18_io_out)
  );
  MyCounter r_count_19 ( // @[SWChisel.scala 171:41]
    .clock(r_count_19_clock),
    .reset(r_count_19_reset),
    .io_en(r_count_19_io_en),
    .io_out(r_count_19_io_out)
  );
  MyCounter r_count_20 ( // @[SWChisel.scala 171:41]
    .clock(r_count_20_clock),
    .reset(r_count_20_reset),
    .io_en(r_count_20_io_en),
    .io_out(r_count_20_io_out)
  );
  MyCounter r_count_21 ( // @[SWChisel.scala 171:41]
    .clock(r_count_21_clock),
    .reset(r_count_21_reset),
    .io_en(r_count_21_io_en),
    .io_out(r_count_21_io_out)
  );
  MyCounter r_count_22 ( // @[SWChisel.scala 171:41]
    .clock(r_count_22_clock),
    .reset(r_count_22_reset),
    .io_en(r_count_22_io_en),
    .io_out(r_count_22_io_out)
  );
  MyCounter r_count_23 ( // @[SWChisel.scala 171:41]
    .clock(r_count_23_clock),
    .reset(r_count_23_reset),
    .io_en(r_count_23_io_en),
    .io_out(r_count_23_io_out)
  );
  MyCounter r_count_24 ( // @[SWChisel.scala 171:41]
    .clock(r_count_24_clock),
    .reset(r_count_24_reset),
    .io_en(r_count_24_io_en),
    .io_out(r_count_24_io_out)
  );
  MyCounter r_count_25 ( // @[SWChisel.scala 171:41]
    .clock(r_count_25_clock),
    .reset(r_count_25_reset),
    .io_en(r_count_25_io_en),
    .io_out(r_count_25_io_out)
  );
  MyCounter r_count_26 ( // @[SWChisel.scala 171:41]
    .clock(r_count_26_clock),
    .reset(r_count_26_reset),
    .io_en(r_count_26_io_en),
    .io_out(r_count_26_io_out)
  );
  MyCounter r_count_27 ( // @[SWChisel.scala 171:41]
    .clock(r_count_27_clock),
    .reset(r_count_27_reset),
    .io_en(r_count_27_io_en),
    .io_out(r_count_27_io_out)
  );
  MyCounter r_count_28 ( // @[SWChisel.scala 171:41]
    .clock(r_count_28_clock),
    .reset(r_count_28_reset),
    .io_en(r_count_28_io_en),
    .io_out(r_count_28_io_out)
  );
  MyCounter r_count_29 ( // @[SWChisel.scala 171:41]
    .clock(r_count_29_clock),
    .reset(r_count_29_reset),
    .io_en(r_count_29_io_en),
    .io_out(r_count_29_io_out)
  );
  MyCounter r_count_30 ( // @[SWChisel.scala 171:41]
    .clock(r_count_30_clock),
    .reset(r_count_30_reset),
    .io_en(r_count_30_io_en),
    .io_out(r_count_30_io_out)
  );
  MyCounter r_count_31 ( // @[SWChisel.scala 171:41]
    .clock(r_count_31_clock),
    .reset(r_count_31_reset),
    .io_en(r_count_31_io_en),
    .io_out(r_count_31_io_out)
  );
  MyCounter r_count_32 ( // @[SWChisel.scala 171:41]
    .clock(r_count_32_clock),
    .reset(r_count_32_reset),
    .io_en(r_count_32_io_en),
    .io_out(r_count_32_io_out)
  );
  MyCounter r_count_33 ( // @[SWChisel.scala 171:41]
    .clock(r_count_33_clock),
    .reset(r_count_33_reset),
    .io_en(r_count_33_io_en),
    .io_out(r_count_33_io_out)
  );
  MyCounter r_count_34 ( // @[SWChisel.scala 171:41]
    .clock(r_count_34_clock),
    .reset(r_count_34_reset),
    .io_en(r_count_34_io_en),
    .io_out(r_count_34_io_out)
  );
  MyCounter r_count_35 ( // @[SWChisel.scala 171:41]
    .clock(r_count_35_clock),
    .reset(r_count_35_reset),
    .io_en(r_count_35_io_en),
    .io_out(r_count_35_io_out)
  );
  MyCounter r_count_36 ( // @[SWChisel.scala 171:41]
    .clock(r_count_36_clock),
    .reset(r_count_36_reset),
    .io_en(r_count_36_io_en),
    .io_out(r_count_36_io_out)
  );
  MyCounter r_count_37 ( // @[SWChisel.scala 171:41]
    .clock(r_count_37_clock),
    .reset(r_count_37_reset),
    .io_en(r_count_37_io_en),
    .io_out(r_count_37_io_out)
  );
  MyCounter r_count_38 ( // @[SWChisel.scala 171:41]
    .clock(r_count_38_clock),
    .reset(r_count_38_reset),
    .io_en(r_count_38_io_en),
    .io_out(r_count_38_io_out)
  );
  MyCounter r_count_39 ( // @[SWChisel.scala 171:41]
    .clock(r_count_39_clock),
    .reset(r_count_39_reset),
    .io_en(r_count_39_io_en),
    .io_out(r_count_39_io_out)
  );
  MyCounter r_count_40 ( // @[SWChisel.scala 171:41]
    .clock(r_count_40_clock),
    .reset(r_count_40_reset),
    .io_en(r_count_40_io_en),
    .io_out(r_count_40_io_out)
  );
  MyCounter r_count_41 ( // @[SWChisel.scala 171:41]
    .clock(r_count_41_clock),
    .reset(r_count_41_reset),
    .io_en(r_count_41_io_en),
    .io_out(r_count_41_io_out)
  );
  MyCounter r_count_42 ( // @[SWChisel.scala 171:41]
    .clock(r_count_42_clock),
    .reset(r_count_42_reset),
    .io_en(r_count_42_io_en),
    .io_out(r_count_42_io_out)
  );
  MyCounter r_count_43 ( // @[SWChisel.scala 171:41]
    .clock(r_count_43_clock),
    .reset(r_count_43_reset),
    .io_en(r_count_43_io_en),
    .io_out(r_count_43_io_out)
  );
  MyCounter r_count_44 ( // @[SWChisel.scala 171:41]
    .clock(r_count_44_clock),
    .reset(r_count_44_reset),
    .io_en(r_count_44_io_en),
    .io_out(r_count_44_io_out)
  );
  MyCounter r_count_45 ( // @[SWChisel.scala 171:41]
    .clock(r_count_45_clock),
    .reset(r_count_45_reset),
    .io_en(r_count_45_io_en),
    .io_out(r_count_45_io_out)
  );
  MyCounter r_count_46 ( // @[SWChisel.scala 171:41]
    .clock(r_count_46_clock),
    .reset(r_count_46_reset),
    .io_en(r_count_46_io_en),
    .io_out(r_count_46_io_out)
  );
  MyCounter r_count_47 ( // @[SWChisel.scala 171:41]
    .clock(r_count_47_clock),
    .reset(r_count_47_reset),
    .io_en(r_count_47_io_en),
    .io_out(r_count_47_io_out)
  );
  MyCounter r_count_48 ( // @[SWChisel.scala 171:41]
    .clock(r_count_48_clock),
    .reset(r_count_48_reset),
    .io_en(r_count_48_io_en),
    .io_out(r_count_48_io_out)
  );
  MyCounter r_count_49 ( // @[SWChisel.scala 171:41]
    .clock(r_count_49_clock),
    .reset(r_count_49_reset),
    .io_en(r_count_49_io_en),
    .io_out(r_count_49_io_out)
  );
  MyCounter r_count_50 ( // @[SWChisel.scala 171:41]
    .clock(r_count_50_clock),
    .reset(r_count_50_reset),
    .io_en(r_count_50_io_en),
    .io_out(r_count_50_io_out)
  );
  MyCounter r_count_51 ( // @[SWChisel.scala 171:41]
    .clock(r_count_51_clock),
    .reset(r_count_51_reset),
    .io_en(r_count_51_io_en),
    .io_out(r_count_51_io_out)
  );
  MyCounter r_count_52 ( // @[SWChisel.scala 171:41]
    .clock(r_count_52_clock),
    .reset(r_count_52_reset),
    .io_en(r_count_52_io_en),
    .io_out(r_count_52_io_out)
  );
  MyCounter r_count_53 ( // @[SWChisel.scala 171:41]
    .clock(r_count_53_clock),
    .reset(r_count_53_reset),
    .io_en(r_count_53_io_en),
    .io_out(r_count_53_io_out)
  );
  MyCounter r_count_54 ( // @[SWChisel.scala 171:41]
    .clock(r_count_54_clock),
    .reset(r_count_54_reset),
    .io_en(r_count_54_io_en),
    .io_out(r_count_54_io_out)
  );
  MyCounter r_count_55 ( // @[SWChisel.scala 171:41]
    .clock(r_count_55_clock),
    .reset(r_count_55_reset),
    .io_en(r_count_55_io_en),
    .io_out(r_count_55_io_out)
  );
  MyCounter r_count_56 ( // @[SWChisel.scala 171:41]
    .clock(r_count_56_clock),
    .reset(r_count_56_reset),
    .io_en(r_count_56_io_en),
    .io_out(r_count_56_io_out)
  );
  MyCounter r_count_57 ( // @[SWChisel.scala 171:41]
    .clock(r_count_57_clock),
    .reset(r_count_57_reset),
    .io_en(r_count_57_io_en),
    .io_out(r_count_57_io_out)
  );
  MyCounter r_count_58 ( // @[SWChisel.scala 171:41]
    .clock(r_count_58_clock),
    .reset(r_count_58_reset),
    .io_en(r_count_58_io_en),
    .io_out(r_count_58_io_out)
  );
  MyCounter r_count_59 ( // @[SWChisel.scala 171:41]
    .clock(r_count_59_clock),
    .reset(r_count_59_reset),
    .io_en(r_count_59_io_en),
    .io_out(r_count_59_io_out)
  );
  MAX max ( // @[SWChisel.scala 174:19]
    .clock(max_clock),
    .reset(max_reset),
    .io_start(max_io_start),
    .io_in(max_io_in),
    .io_done(max_io_done),
    .io_out(max_io_out)
  );
  assign io_result = max_io_out; // @[SWChisel.scala 181:13]
  assign io_done = max_io_done; // @[SWChisel.scala 182:11]
  assign array_0_io_q = io_q_0_b; // @[SWChisel.scala 220:19]
  assign array_0_io_r = 9'h18f == r_count_0_io_out ? io_r_399_b : _GEN_578; // @[SWChisel.scala 221:{19,19}]
  assign array_0_io_e_i = E_0; // @[SWChisel.scala 196:21]
  assign array_0_io_f_i = 16'sh0; // @[SWChisel.scala 198:21]
  assign array_0_io_ve_i = V1_1; // @[SWChisel.scala 197:22]
  assign array_0_io_vf_i = V1_0; // @[SWChisel.scala 199:22]
  assign array_0_io_vv_i = V2_0; // @[SWChisel.scala 200:22]
  assign array_1_io_q = io_q_1_b; // @[SWChisel.scala 220:19]
  assign array_1_io_r = 9'h18f == r_count_1_io_out ? io_r_399_b : _GEN_978; // @[SWChisel.scala 221:{19,19}]
  assign array_1_io_e_i = E_1; // @[SWChisel.scala 196:21]
  assign array_1_io_f_i = F_1; // @[SWChisel.scala 198:21]
  assign array_1_io_ve_i = V1_2; // @[SWChisel.scala 197:22]
  assign array_1_io_vf_i = V1_1; // @[SWChisel.scala 199:22]
  assign array_1_io_vv_i = V2_1; // @[SWChisel.scala 200:22]
  assign array_2_io_q = io_q_2_b; // @[SWChisel.scala 220:19]
  assign array_2_io_r = 9'h18f == r_count_2_io_out ? io_r_399_b : _GEN_1378; // @[SWChisel.scala 221:{19,19}]
  assign array_2_io_e_i = E_2; // @[SWChisel.scala 196:21]
  assign array_2_io_f_i = F_2; // @[SWChisel.scala 198:21]
  assign array_2_io_ve_i = V1_3; // @[SWChisel.scala 197:22]
  assign array_2_io_vf_i = V1_2; // @[SWChisel.scala 199:22]
  assign array_2_io_vv_i = V2_2; // @[SWChisel.scala 200:22]
  assign array_3_io_q = io_q_3_b; // @[SWChisel.scala 220:19]
  assign array_3_io_r = 9'h18f == r_count_3_io_out ? io_r_399_b : _GEN_1778; // @[SWChisel.scala 221:{19,19}]
  assign array_3_io_e_i = E_3; // @[SWChisel.scala 196:21]
  assign array_3_io_f_i = F_3; // @[SWChisel.scala 198:21]
  assign array_3_io_ve_i = V1_4; // @[SWChisel.scala 197:22]
  assign array_3_io_vf_i = V1_3; // @[SWChisel.scala 199:22]
  assign array_3_io_vv_i = V2_3; // @[SWChisel.scala 200:22]
  assign array_4_io_q = io_q_4_b; // @[SWChisel.scala 220:19]
  assign array_4_io_r = 9'h18f == r_count_4_io_out ? io_r_399_b : _GEN_2178; // @[SWChisel.scala 221:{19,19}]
  assign array_4_io_e_i = E_4; // @[SWChisel.scala 196:21]
  assign array_4_io_f_i = F_4; // @[SWChisel.scala 198:21]
  assign array_4_io_ve_i = V1_5; // @[SWChisel.scala 197:22]
  assign array_4_io_vf_i = V1_4; // @[SWChisel.scala 199:22]
  assign array_4_io_vv_i = V2_4; // @[SWChisel.scala 200:22]
  assign array_5_io_q = io_q_5_b; // @[SWChisel.scala 220:19]
  assign array_5_io_r = 9'h18f == r_count_5_io_out ? io_r_399_b : _GEN_2578; // @[SWChisel.scala 221:{19,19}]
  assign array_5_io_e_i = E_5; // @[SWChisel.scala 196:21]
  assign array_5_io_f_i = F_5; // @[SWChisel.scala 198:21]
  assign array_5_io_ve_i = V1_6; // @[SWChisel.scala 197:22]
  assign array_5_io_vf_i = V1_5; // @[SWChisel.scala 199:22]
  assign array_5_io_vv_i = V2_5; // @[SWChisel.scala 200:22]
  assign array_6_io_q = io_q_6_b; // @[SWChisel.scala 220:19]
  assign array_6_io_r = 9'h18f == r_count_6_io_out ? io_r_399_b : _GEN_2978; // @[SWChisel.scala 221:{19,19}]
  assign array_6_io_e_i = E_6; // @[SWChisel.scala 196:21]
  assign array_6_io_f_i = F_6; // @[SWChisel.scala 198:21]
  assign array_6_io_ve_i = V1_7; // @[SWChisel.scala 197:22]
  assign array_6_io_vf_i = V1_6; // @[SWChisel.scala 199:22]
  assign array_6_io_vv_i = V2_6; // @[SWChisel.scala 200:22]
  assign array_7_io_q = io_q_7_b; // @[SWChisel.scala 220:19]
  assign array_7_io_r = 9'h18f == r_count_7_io_out ? io_r_399_b : _GEN_3378; // @[SWChisel.scala 221:{19,19}]
  assign array_7_io_e_i = E_7; // @[SWChisel.scala 196:21]
  assign array_7_io_f_i = F_7; // @[SWChisel.scala 198:21]
  assign array_7_io_ve_i = V1_8; // @[SWChisel.scala 197:22]
  assign array_7_io_vf_i = V1_7; // @[SWChisel.scala 199:22]
  assign array_7_io_vv_i = V2_7; // @[SWChisel.scala 200:22]
  assign array_8_io_q = io_q_8_b; // @[SWChisel.scala 220:19]
  assign array_8_io_r = 9'h18f == r_count_8_io_out ? io_r_399_b : _GEN_3778; // @[SWChisel.scala 221:{19,19}]
  assign array_8_io_e_i = E_8; // @[SWChisel.scala 196:21]
  assign array_8_io_f_i = F_8; // @[SWChisel.scala 198:21]
  assign array_8_io_ve_i = V1_9; // @[SWChisel.scala 197:22]
  assign array_8_io_vf_i = V1_8; // @[SWChisel.scala 199:22]
  assign array_8_io_vv_i = V2_8; // @[SWChisel.scala 200:22]
  assign array_9_io_q = io_q_9_b; // @[SWChisel.scala 220:19]
  assign array_9_io_r = 9'h18f == r_count_9_io_out ? io_r_399_b : _GEN_4178; // @[SWChisel.scala 221:{19,19}]
  assign array_9_io_e_i = E_9; // @[SWChisel.scala 196:21]
  assign array_9_io_f_i = F_9; // @[SWChisel.scala 198:21]
  assign array_9_io_ve_i = V1_10; // @[SWChisel.scala 197:22]
  assign array_9_io_vf_i = V1_9; // @[SWChisel.scala 199:22]
  assign array_9_io_vv_i = V2_9; // @[SWChisel.scala 200:22]
  assign array_10_io_q = io_q_10_b; // @[SWChisel.scala 220:19]
  assign array_10_io_r = 9'h18f == r_count_10_io_out ? io_r_399_b : _GEN_4578; // @[SWChisel.scala 221:{19,19}]
  assign array_10_io_e_i = E_10; // @[SWChisel.scala 196:21]
  assign array_10_io_f_i = F_10; // @[SWChisel.scala 198:21]
  assign array_10_io_ve_i = V1_11; // @[SWChisel.scala 197:22]
  assign array_10_io_vf_i = V1_10; // @[SWChisel.scala 199:22]
  assign array_10_io_vv_i = V2_10; // @[SWChisel.scala 200:22]
  assign array_11_io_q = io_q_11_b; // @[SWChisel.scala 220:19]
  assign array_11_io_r = 9'h18f == r_count_11_io_out ? io_r_399_b : _GEN_4978; // @[SWChisel.scala 221:{19,19}]
  assign array_11_io_e_i = E_11; // @[SWChisel.scala 196:21]
  assign array_11_io_f_i = F_11; // @[SWChisel.scala 198:21]
  assign array_11_io_ve_i = V1_12; // @[SWChisel.scala 197:22]
  assign array_11_io_vf_i = V1_11; // @[SWChisel.scala 199:22]
  assign array_11_io_vv_i = V2_11; // @[SWChisel.scala 200:22]
  assign array_12_io_q = io_q_12_b; // @[SWChisel.scala 220:19]
  assign array_12_io_r = 9'h18f == r_count_12_io_out ? io_r_399_b : _GEN_5378; // @[SWChisel.scala 221:{19,19}]
  assign array_12_io_e_i = E_12; // @[SWChisel.scala 196:21]
  assign array_12_io_f_i = F_12; // @[SWChisel.scala 198:21]
  assign array_12_io_ve_i = V1_13; // @[SWChisel.scala 197:22]
  assign array_12_io_vf_i = V1_12; // @[SWChisel.scala 199:22]
  assign array_12_io_vv_i = V2_12; // @[SWChisel.scala 200:22]
  assign array_13_io_q = io_q_13_b; // @[SWChisel.scala 220:19]
  assign array_13_io_r = 9'h18f == r_count_13_io_out ? io_r_399_b : _GEN_5778; // @[SWChisel.scala 221:{19,19}]
  assign array_13_io_e_i = E_13; // @[SWChisel.scala 196:21]
  assign array_13_io_f_i = F_13; // @[SWChisel.scala 198:21]
  assign array_13_io_ve_i = V1_14; // @[SWChisel.scala 197:22]
  assign array_13_io_vf_i = V1_13; // @[SWChisel.scala 199:22]
  assign array_13_io_vv_i = V2_13; // @[SWChisel.scala 200:22]
  assign array_14_io_q = io_q_14_b; // @[SWChisel.scala 220:19]
  assign array_14_io_r = 9'h18f == r_count_14_io_out ? io_r_399_b : _GEN_6178; // @[SWChisel.scala 221:{19,19}]
  assign array_14_io_e_i = E_14; // @[SWChisel.scala 196:21]
  assign array_14_io_f_i = F_14; // @[SWChisel.scala 198:21]
  assign array_14_io_ve_i = V1_15; // @[SWChisel.scala 197:22]
  assign array_14_io_vf_i = V1_14; // @[SWChisel.scala 199:22]
  assign array_14_io_vv_i = V2_14; // @[SWChisel.scala 200:22]
  assign array_15_io_q = io_q_15_b; // @[SWChisel.scala 220:19]
  assign array_15_io_r = 9'h18f == r_count_15_io_out ? io_r_399_b : _GEN_6578; // @[SWChisel.scala 221:{19,19}]
  assign array_15_io_e_i = E_15; // @[SWChisel.scala 196:21]
  assign array_15_io_f_i = F_15; // @[SWChisel.scala 198:21]
  assign array_15_io_ve_i = V1_16; // @[SWChisel.scala 197:22]
  assign array_15_io_vf_i = V1_15; // @[SWChisel.scala 199:22]
  assign array_15_io_vv_i = V2_15; // @[SWChisel.scala 200:22]
  assign array_16_io_q = io_q_16_b; // @[SWChisel.scala 220:19]
  assign array_16_io_r = 9'h18f == r_count_16_io_out ? io_r_399_b : _GEN_6978; // @[SWChisel.scala 221:{19,19}]
  assign array_16_io_e_i = E_16; // @[SWChisel.scala 196:21]
  assign array_16_io_f_i = F_16; // @[SWChisel.scala 198:21]
  assign array_16_io_ve_i = V1_17; // @[SWChisel.scala 197:22]
  assign array_16_io_vf_i = V1_16; // @[SWChisel.scala 199:22]
  assign array_16_io_vv_i = V2_16; // @[SWChisel.scala 200:22]
  assign array_17_io_q = io_q_17_b; // @[SWChisel.scala 220:19]
  assign array_17_io_r = 9'h18f == r_count_17_io_out ? io_r_399_b : _GEN_7378; // @[SWChisel.scala 221:{19,19}]
  assign array_17_io_e_i = E_17; // @[SWChisel.scala 196:21]
  assign array_17_io_f_i = F_17; // @[SWChisel.scala 198:21]
  assign array_17_io_ve_i = V1_18; // @[SWChisel.scala 197:22]
  assign array_17_io_vf_i = V1_17; // @[SWChisel.scala 199:22]
  assign array_17_io_vv_i = V2_17; // @[SWChisel.scala 200:22]
  assign array_18_io_q = io_q_18_b; // @[SWChisel.scala 220:19]
  assign array_18_io_r = 9'h18f == r_count_18_io_out ? io_r_399_b : _GEN_7778; // @[SWChisel.scala 221:{19,19}]
  assign array_18_io_e_i = E_18; // @[SWChisel.scala 196:21]
  assign array_18_io_f_i = F_18; // @[SWChisel.scala 198:21]
  assign array_18_io_ve_i = V1_19; // @[SWChisel.scala 197:22]
  assign array_18_io_vf_i = V1_18; // @[SWChisel.scala 199:22]
  assign array_18_io_vv_i = V2_18; // @[SWChisel.scala 200:22]
  assign array_19_io_q = io_q_19_b; // @[SWChisel.scala 220:19]
  assign array_19_io_r = 9'h18f == r_count_19_io_out ? io_r_399_b : _GEN_8178; // @[SWChisel.scala 221:{19,19}]
  assign array_19_io_e_i = E_19; // @[SWChisel.scala 196:21]
  assign array_19_io_f_i = F_19; // @[SWChisel.scala 198:21]
  assign array_19_io_ve_i = V1_20; // @[SWChisel.scala 197:22]
  assign array_19_io_vf_i = V1_19; // @[SWChisel.scala 199:22]
  assign array_19_io_vv_i = V2_19; // @[SWChisel.scala 200:22]
  assign array_20_io_q = io_q_20_b; // @[SWChisel.scala 220:19]
  assign array_20_io_r = 9'h18f == r_count_20_io_out ? io_r_399_b : _GEN_8578; // @[SWChisel.scala 221:{19,19}]
  assign array_20_io_e_i = E_20; // @[SWChisel.scala 196:21]
  assign array_20_io_f_i = F_20; // @[SWChisel.scala 198:21]
  assign array_20_io_ve_i = V1_21; // @[SWChisel.scala 197:22]
  assign array_20_io_vf_i = V1_20; // @[SWChisel.scala 199:22]
  assign array_20_io_vv_i = V2_20; // @[SWChisel.scala 200:22]
  assign array_21_io_q = io_q_21_b; // @[SWChisel.scala 220:19]
  assign array_21_io_r = 9'h18f == r_count_21_io_out ? io_r_399_b : _GEN_8978; // @[SWChisel.scala 221:{19,19}]
  assign array_21_io_e_i = E_21; // @[SWChisel.scala 196:21]
  assign array_21_io_f_i = F_21; // @[SWChisel.scala 198:21]
  assign array_21_io_ve_i = V1_22; // @[SWChisel.scala 197:22]
  assign array_21_io_vf_i = V1_21; // @[SWChisel.scala 199:22]
  assign array_21_io_vv_i = V2_21; // @[SWChisel.scala 200:22]
  assign array_22_io_q = io_q_22_b; // @[SWChisel.scala 220:19]
  assign array_22_io_r = 9'h18f == r_count_22_io_out ? io_r_399_b : _GEN_9378; // @[SWChisel.scala 221:{19,19}]
  assign array_22_io_e_i = E_22; // @[SWChisel.scala 196:21]
  assign array_22_io_f_i = F_22; // @[SWChisel.scala 198:21]
  assign array_22_io_ve_i = V1_23; // @[SWChisel.scala 197:22]
  assign array_22_io_vf_i = V1_22; // @[SWChisel.scala 199:22]
  assign array_22_io_vv_i = V2_22; // @[SWChisel.scala 200:22]
  assign array_23_io_q = io_q_23_b; // @[SWChisel.scala 220:19]
  assign array_23_io_r = 9'h18f == r_count_23_io_out ? io_r_399_b : _GEN_9778; // @[SWChisel.scala 221:{19,19}]
  assign array_23_io_e_i = E_23; // @[SWChisel.scala 196:21]
  assign array_23_io_f_i = F_23; // @[SWChisel.scala 198:21]
  assign array_23_io_ve_i = V1_24; // @[SWChisel.scala 197:22]
  assign array_23_io_vf_i = V1_23; // @[SWChisel.scala 199:22]
  assign array_23_io_vv_i = V2_23; // @[SWChisel.scala 200:22]
  assign array_24_io_q = io_q_24_b; // @[SWChisel.scala 220:19]
  assign array_24_io_r = 9'h18f == r_count_24_io_out ? io_r_399_b : _GEN_10178; // @[SWChisel.scala 221:{19,19}]
  assign array_24_io_e_i = E_24; // @[SWChisel.scala 196:21]
  assign array_24_io_f_i = F_24; // @[SWChisel.scala 198:21]
  assign array_24_io_ve_i = V1_25; // @[SWChisel.scala 197:22]
  assign array_24_io_vf_i = V1_24; // @[SWChisel.scala 199:22]
  assign array_24_io_vv_i = V2_24; // @[SWChisel.scala 200:22]
  assign array_25_io_q = io_q_25_b; // @[SWChisel.scala 220:19]
  assign array_25_io_r = 9'h18f == r_count_25_io_out ? io_r_399_b : _GEN_10578; // @[SWChisel.scala 221:{19,19}]
  assign array_25_io_e_i = E_25; // @[SWChisel.scala 196:21]
  assign array_25_io_f_i = F_25; // @[SWChisel.scala 198:21]
  assign array_25_io_ve_i = V1_26; // @[SWChisel.scala 197:22]
  assign array_25_io_vf_i = V1_25; // @[SWChisel.scala 199:22]
  assign array_25_io_vv_i = V2_25; // @[SWChisel.scala 200:22]
  assign array_26_io_q = io_q_26_b; // @[SWChisel.scala 220:19]
  assign array_26_io_r = 9'h18f == r_count_26_io_out ? io_r_399_b : _GEN_10978; // @[SWChisel.scala 221:{19,19}]
  assign array_26_io_e_i = E_26; // @[SWChisel.scala 196:21]
  assign array_26_io_f_i = F_26; // @[SWChisel.scala 198:21]
  assign array_26_io_ve_i = V1_27; // @[SWChisel.scala 197:22]
  assign array_26_io_vf_i = V1_26; // @[SWChisel.scala 199:22]
  assign array_26_io_vv_i = V2_26; // @[SWChisel.scala 200:22]
  assign array_27_io_q = io_q_27_b; // @[SWChisel.scala 220:19]
  assign array_27_io_r = 9'h18f == r_count_27_io_out ? io_r_399_b : _GEN_11378; // @[SWChisel.scala 221:{19,19}]
  assign array_27_io_e_i = E_27; // @[SWChisel.scala 196:21]
  assign array_27_io_f_i = F_27; // @[SWChisel.scala 198:21]
  assign array_27_io_ve_i = V1_28; // @[SWChisel.scala 197:22]
  assign array_27_io_vf_i = V1_27; // @[SWChisel.scala 199:22]
  assign array_27_io_vv_i = V2_27; // @[SWChisel.scala 200:22]
  assign array_28_io_q = io_q_28_b; // @[SWChisel.scala 220:19]
  assign array_28_io_r = 9'h18f == r_count_28_io_out ? io_r_399_b : _GEN_11778; // @[SWChisel.scala 221:{19,19}]
  assign array_28_io_e_i = E_28; // @[SWChisel.scala 196:21]
  assign array_28_io_f_i = F_28; // @[SWChisel.scala 198:21]
  assign array_28_io_ve_i = V1_29; // @[SWChisel.scala 197:22]
  assign array_28_io_vf_i = V1_28; // @[SWChisel.scala 199:22]
  assign array_28_io_vv_i = V2_28; // @[SWChisel.scala 200:22]
  assign array_29_io_q = io_q_29_b; // @[SWChisel.scala 220:19]
  assign array_29_io_r = 9'h18f == r_count_29_io_out ? io_r_399_b : _GEN_12178; // @[SWChisel.scala 221:{19,19}]
  assign array_29_io_e_i = E_29; // @[SWChisel.scala 196:21]
  assign array_29_io_f_i = F_29; // @[SWChisel.scala 198:21]
  assign array_29_io_ve_i = V1_30; // @[SWChisel.scala 197:22]
  assign array_29_io_vf_i = V1_29; // @[SWChisel.scala 199:22]
  assign array_29_io_vv_i = V2_29; // @[SWChisel.scala 200:22]
  assign array_30_io_q = io_q_30_b; // @[SWChisel.scala 220:19]
  assign array_30_io_r = 9'h18f == r_count_30_io_out ? io_r_399_b : _GEN_12578; // @[SWChisel.scala 221:{19,19}]
  assign array_30_io_e_i = E_30; // @[SWChisel.scala 196:21]
  assign array_30_io_f_i = F_30; // @[SWChisel.scala 198:21]
  assign array_30_io_ve_i = V1_31; // @[SWChisel.scala 197:22]
  assign array_30_io_vf_i = V1_30; // @[SWChisel.scala 199:22]
  assign array_30_io_vv_i = V2_30; // @[SWChisel.scala 200:22]
  assign array_31_io_q = io_q_31_b; // @[SWChisel.scala 220:19]
  assign array_31_io_r = 9'h18f == r_count_31_io_out ? io_r_399_b : _GEN_12978; // @[SWChisel.scala 221:{19,19}]
  assign array_31_io_e_i = E_31; // @[SWChisel.scala 196:21]
  assign array_31_io_f_i = F_31; // @[SWChisel.scala 198:21]
  assign array_31_io_ve_i = V1_32; // @[SWChisel.scala 197:22]
  assign array_31_io_vf_i = V1_31; // @[SWChisel.scala 199:22]
  assign array_31_io_vv_i = V2_31; // @[SWChisel.scala 200:22]
  assign array_32_io_q = io_q_32_b; // @[SWChisel.scala 220:19]
  assign array_32_io_r = 9'h18f == r_count_32_io_out ? io_r_399_b : _GEN_13378; // @[SWChisel.scala 221:{19,19}]
  assign array_32_io_e_i = E_32; // @[SWChisel.scala 196:21]
  assign array_32_io_f_i = F_32; // @[SWChisel.scala 198:21]
  assign array_32_io_ve_i = V1_33; // @[SWChisel.scala 197:22]
  assign array_32_io_vf_i = V1_32; // @[SWChisel.scala 199:22]
  assign array_32_io_vv_i = V2_32; // @[SWChisel.scala 200:22]
  assign array_33_io_q = io_q_33_b; // @[SWChisel.scala 220:19]
  assign array_33_io_r = 9'h18f == r_count_33_io_out ? io_r_399_b : _GEN_13778; // @[SWChisel.scala 221:{19,19}]
  assign array_33_io_e_i = E_33; // @[SWChisel.scala 196:21]
  assign array_33_io_f_i = F_33; // @[SWChisel.scala 198:21]
  assign array_33_io_ve_i = V1_34; // @[SWChisel.scala 197:22]
  assign array_33_io_vf_i = V1_33; // @[SWChisel.scala 199:22]
  assign array_33_io_vv_i = V2_33; // @[SWChisel.scala 200:22]
  assign array_34_io_q = io_q_34_b; // @[SWChisel.scala 220:19]
  assign array_34_io_r = 9'h18f == r_count_34_io_out ? io_r_399_b : _GEN_14178; // @[SWChisel.scala 221:{19,19}]
  assign array_34_io_e_i = E_34; // @[SWChisel.scala 196:21]
  assign array_34_io_f_i = F_34; // @[SWChisel.scala 198:21]
  assign array_34_io_ve_i = V1_35; // @[SWChisel.scala 197:22]
  assign array_34_io_vf_i = V1_34; // @[SWChisel.scala 199:22]
  assign array_34_io_vv_i = V2_34; // @[SWChisel.scala 200:22]
  assign array_35_io_q = io_q_35_b; // @[SWChisel.scala 220:19]
  assign array_35_io_r = 9'h18f == r_count_35_io_out ? io_r_399_b : _GEN_14578; // @[SWChisel.scala 221:{19,19}]
  assign array_35_io_e_i = E_35; // @[SWChisel.scala 196:21]
  assign array_35_io_f_i = F_35; // @[SWChisel.scala 198:21]
  assign array_35_io_ve_i = V1_36; // @[SWChisel.scala 197:22]
  assign array_35_io_vf_i = V1_35; // @[SWChisel.scala 199:22]
  assign array_35_io_vv_i = V2_35; // @[SWChisel.scala 200:22]
  assign array_36_io_q = io_q_36_b; // @[SWChisel.scala 220:19]
  assign array_36_io_r = 9'h18f == r_count_36_io_out ? io_r_399_b : _GEN_14978; // @[SWChisel.scala 221:{19,19}]
  assign array_36_io_e_i = E_36; // @[SWChisel.scala 196:21]
  assign array_36_io_f_i = F_36; // @[SWChisel.scala 198:21]
  assign array_36_io_ve_i = V1_37; // @[SWChisel.scala 197:22]
  assign array_36_io_vf_i = V1_36; // @[SWChisel.scala 199:22]
  assign array_36_io_vv_i = V2_36; // @[SWChisel.scala 200:22]
  assign array_37_io_q = io_q_37_b; // @[SWChisel.scala 220:19]
  assign array_37_io_r = 9'h18f == r_count_37_io_out ? io_r_399_b : _GEN_15378; // @[SWChisel.scala 221:{19,19}]
  assign array_37_io_e_i = E_37; // @[SWChisel.scala 196:21]
  assign array_37_io_f_i = F_37; // @[SWChisel.scala 198:21]
  assign array_37_io_ve_i = V1_38; // @[SWChisel.scala 197:22]
  assign array_37_io_vf_i = V1_37; // @[SWChisel.scala 199:22]
  assign array_37_io_vv_i = V2_37; // @[SWChisel.scala 200:22]
  assign array_38_io_q = io_q_38_b; // @[SWChisel.scala 220:19]
  assign array_38_io_r = 9'h18f == r_count_38_io_out ? io_r_399_b : _GEN_15778; // @[SWChisel.scala 221:{19,19}]
  assign array_38_io_e_i = E_38; // @[SWChisel.scala 196:21]
  assign array_38_io_f_i = F_38; // @[SWChisel.scala 198:21]
  assign array_38_io_ve_i = V1_39; // @[SWChisel.scala 197:22]
  assign array_38_io_vf_i = V1_38; // @[SWChisel.scala 199:22]
  assign array_38_io_vv_i = V2_38; // @[SWChisel.scala 200:22]
  assign array_39_io_q = io_q_39_b; // @[SWChisel.scala 220:19]
  assign array_39_io_r = 9'h18f == r_count_39_io_out ? io_r_399_b : _GEN_16178; // @[SWChisel.scala 221:{19,19}]
  assign array_39_io_e_i = E_39; // @[SWChisel.scala 196:21]
  assign array_39_io_f_i = F_39; // @[SWChisel.scala 198:21]
  assign array_39_io_ve_i = V1_40; // @[SWChisel.scala 197:22]
  assign array_39_io_vf_i = V1_39; // @[SWChisel.scala 199:22]
  assign array_39_io_vv_i = V2_39; // @[SWChisel.scala 200:22]
  assign array_40_io_q = io_q_40_b; // @[SWChisel.scala 220:19]
  assign array_40_io_r = 9'h18f == r_count_40_io_out ? io_r_399_b : _GEN_16578; // @[SWChisel.scala 221:{19,19}]
  assign array_40_io_e_i = E_40; // @[SWChisel.scala 196:21]
  assign array_40_io_f_i = F_40; // @[SWChisel.scala 198:21]
  assign array_40_io_ve_i = V1_41; // @[SWChisel.scala 197:22]
  assign array_40_io_vf_i = V1_40; // @[SWChisel.scala 199:22]
  assign array_40_io_vv_i = V2_40; // @[SWChisel.scala 200:22]
  assign array_41_io_q = io_q_41_b; // @[SWChisel.scala 220:19]
  assign array_41_io_r = 9'h18f == r_count_41_io_out ? io_r_399_b : _GEN_16978; // @[SWChisel.scala 221:{19,19}]
  assign array_41_io_e_i = E_41; // @[SWChisel.scala 196:21]
  assign array_41_io_f_i = F_41; // @[SWChisel.scala 198:21]
  assign array_41_io_ve_i = V1_42; // @[SWChisel.scala 197:22]
  assign array_41_io_vf_i = V1_41; // @[SWChisel.scala 199:22]
  assign array_41_io_vv_i = V2_41; // @[SWChisel.scala 200:22]
  assign array_42_io_q = io_q_42_b; // @[SWChisel.scala 220:19]
  assign array_42_io_r = 9'h18f == r_count_42_io_out ? io_r_399_b : _GEN_17378; // @[SWChisel.scala 221:{19,19}]
  assign array_42_io_e_i = E_42; // @[SWChisel.scala 196:21]
  assign array_42_io_f_i = F_42; // @[SWChisel.scala 198:21]
  assign array_42_io_ve_i = V1_43; // @[SWChisel.scala 197:22]
  assign array_42_io_vf_i = V1_42; // @[SWChisel.scala 199:22]
  assign array_42_io_vv_i = V2_42; // @[SWChisel.scala 200:22]
  assign array_43_io_q = io_q_43_b; // @[SWChisel.scala 220:19]
  assign array_43_io_r = 9'h18f == r_count_43_io_out ? io_r_399_b : _GEN_17778; // @[SWChisel.scala 221:{19,19}]
  assign array_43_io_e_i = E_43; // @[SWChisel.scala 196:21]
  assign array_43_io_f_i = F_43; // @[SWChisel.scala 198:21]
  assign array_43_io_ve_i = V1_44; // @[SWChisel.scala 197:22]
  assign array_43_io_vf_i = V1_43; // @[SWChisel.scala 199:22]
  assign array_43_io_vv_i = V2_43; // @[SWChisel.scala 200:22]
  assign array_44_io_q = io_q_44_b; // @[SWChisel.scala 220:19]
  assign array_44_io_r = 9'h18f == r_count_44_io_out ? io_r_399_b : _GEN_18178; // @[SWChisel.scala 221:{19,19}]
  assign array_44_io_e_i = E_44; // @[SWChisel.scala 196:21]
  assign array_44_io_f_i = F_44; // @[SWChisel.scala 198:21]
  assign array_44_io_ve_i = V1_45; // @[SWChisel.scala 197:22]
  assign array_44_io_vf_i = V1_44; // @[SWChisel.scala 199:22]
  assign array_44_io_vv_i = V2_44; // @[SWChisel.scala 200:22]
  assign array_45_io_q = io_q_45_b; // @[SWChisel.scala 220:19]
  assign array_45_io_r = 9'h18f == r_count_45_io_out ? io_r_399_b : _GEN_18578; // @[SWChisel.scala 221:{19,19}]
  assign array_45_io_e_i = E_45; // @[SWChisel.scala 196:21]
  assign array_45_io_f_i = F_45; // @[SWChisel.scala 198:21]
  assign array_45_io_ve_i = V1_46; // @[SWChisel.scala 197:22]
  assign array_45_io_vf_i = V1_45; // @[SWChisel.scala 199:22]
  assign array_45_io_vv_i = V2_45; // @[SWChisel.scala 200:22]
  assign array_46_io_q = io_q_46_b; // @[SWChisel.scala 220:19]
  assign array_46_io_r = 9'h18f == r_count_46_io_out ? io_r_399_b : _GEN_18978; // @[SWChisel.scala 221:{19,19}]
  assign array_46_io_e_i = E_46; // @[SWChisel.scala 196:21]
  assign array_46_io_f_i = F_46; // @[SWChisel.scala 198:21]
  assign array_46_io_ve_i = V1_47; // @[SWChisel.scala 197:22]
  assign array_46_io_vf_i = V1_46; // @[SWChisel.scala 199:22]
  assign array_46_io_vv_i = V2_46; // @[SWChisel.scala 200:22]
  assign array_47_io_q = io_q_47_b; // @[SWChisel.scala 220:19]
  assign array_47_io_r = 9'h18f == r_count_47_io_out ? io_r_399_b : _GEN_19378; // @[SWChisel.scala 221:{19,19}]
  assign array_47_io_e_i = E_47; // @[SWChisel.scala 196:21]
  assign array_47_io_f_i = F_47; // @[SWChisel.scala 198:21]
  assign array_47_io_ve_i = V1_48; // @[SWChisel.scala 197:22]
  assign array_47_io_vf_i = V1_47; // @[SWChisel.scala 199:22]
  assign array_47_io_vv_i = V2_47; // @[SWChisel.scala 200:22]
  assign array_48_io_q = io_q_48_b; // @[SWChisel.scala 220:19]
  assign array_48_io_r = 9'h18f == r_count_48_io_out ? io_r_399_b : _GEN_19778; // @[SWChisel.scala 221:{19,19}]
  assign array_48_io_e_i = E_48; // @[SWChisel.scala 196:21]
  assign array_48_io_f_i = F_48; // @[SWChisel.scala 198:21]
  assign array_48_io_ve_i = V1_49; // @[SWChisel.scala 197:22]
  assign array_48_io_vf_i = V1_48; // @[SWChisel.scala 199:22]
  assign array_48_io_vv_i = V2_48; // @[SWChisel.scala 200:22]
  assign array_49_io_q = io_q_49_b; // @[SWChisel.scala 220:19]
  assign array_49_io_r = 9'h18f == r_count_49_io_out ? io_r_399_b : _GEN_20178; // @[SWChisel.scala 221:{19,19}]
  assign array_49_io_e_i = E_49; // @[SWChisel.scala 196:21]
  assign array_49_io_f_i = F_49; // @[SWChisel.scala 198:21]
  assign array_49_io_ve_i = V1_50; // @[SWChisel.scala 197:22]
  assign array_49_io_vf_i = V1_49; // @[SWChisel.scala 199:22]
  assign array_49_io_vv_i = V2_49; // @[SWChisel.scala 200:22]
  assign array_50_io_q = io_q_50_b; // @[SWChisel.scala 220:19]
  assign array_50_io_r = 9'h18f == r_count_50_io_out ? io_r_399_b : _GEN_20578; // @[SWChisel.scala 221:{19,19}]
  assign array_50_io_e_i = E_50; // @[SWChisel.scala 196:21]
  assign array_50_io_f_i = F_50; // @[SWChisel.scala 198:21]
  assign array_50_io_ve_i = V1_51; // @[SWChisel.scala 197:22]
  assign array_50_io_vf_i = V1_50; // @[SWChisel.scala 199:22]
  assign array_50_io_vv_i = V2_50; // @[SWChisel.scala 200:22]
  assign array_51_io_q = io_q_51_b; // @[SWChisel.scala 220:19]
  assign array_51_io_r = 9'h18f == r_count_51_io_out ? io_r_399_b : _GEN_20978; // @[SWChisel.scala 221:{19,19}]
  assign array_51_io_e_i = E_51; // @[SWChisel.scala 196:21]
  assign array_51_io_f_i = F_51; // @[SWChisel.scala 198:21]
  assign array_51_io_ve_i = V1_52; // @[SWChisel.scala 197:22]
  assign array_51_io_vf_i = V1_51; // @[SWChisel.scala 199:22]
  assign array_51_io_vv_i = V2_51; // @[SWChisel.scala 200:22]
  assign array_52_io_q = io_q_52_b; // @[SWChisel.scala 220:19]
  assign array_52_io_r = 9'h18f == r_count_52_io_out ? io_r_399_b : _GEN_21378; // @[SWChisel.scala 221:{19,19}]
  assign array_52_io_e_i = E_52; // @[SWChisel.scala 196:21]
  assign array_52_io_f_i = F_52; // @[SWChisel.scala 198:21]
  assign array_52_io_ve_i = V1_53; // @[SWChisel.scala 197:22]
  assign array_52_io_vf_i = V1_52; // @[SWChisel.scala 199:22]
  assign array_52_io_vv_i = V2_52; // @[SWChisel.scala 200:22]
  assign array_53_io_q = io_q_53_b; // @[SWChisel.scala 220:19]
  assign array_53_io_r = 9'h18f == r_count_53_io_out ? io_r_399_b : _GEN_21778; // @[SWChisel.scala 221:{19,19}]
  assign array_53_io_e_i = E_53; // @[SWChisel.scala 196:21]
  assign array_53_io_f_i = F_53; // @[SWChisel.scala 198:21]
  assign array_53_io_ve_i = V1_54; // @[SWChisel.scala 197:22]
  assign array_53_io_vf_i = V1_53; // @[SWChisel.scala 199:22]
  assign array_53_io_vv_i = V2_53; // @[SWChisel.scala 200:22]
  assign array_54_io_q = io_q_54_b; // @[SWChisel.scala 220:19]
  assign array_54_io_r = 9'h18f == r_count_54_io_out ? io_r_399_b : _GEN_22178; // @[SWChisel.scala 221:{19,19}]
  assign array_54_io_e_i = E_54; // @[SWChisel.scala 196:21]
  assign array_54_io_f_i = F_54; // @[SWChisel.scala 198:21]
  assign array_54_io_ve_i = V1_55; // @[SWChisel.scala 197:22]
  assign array_54_io_vf_i = V1_54; // @[SWChisel.scala 199:22]
  assign array_54_io_vv_i = V2_54; // @[SWChisel.scala 200:22]
  assign array_55_io_q = io_q_55_b; // @[SWChisel.scala 220:19]
  assign array_55_io_r = 9'h18f == r_count_55_io_out ? io_r_399_b : _GEN_22578; // @[SWChisel.scala 221:{19,19}]
  assign array_55_io_e_i = E_55; // @[SWChisel.scala 196:21]
  assign array_55_io_f_i = F_55; // @[SWChisel.scala 198:21]
  assign array_55_io_ve_i = V1_56; // @[SWChisel.scala 197:22]
  assign array_55_io_vf_i = V1_55; // @[SWChisel.scala 199:22]
  assign array_55_io_vv_i = V2_55; // @[SWChisel.scala 200:22]
  assign array_56_io_q = io_q_56_b; // @[SWChisel.scala 220:19]
  assign array_56_io_r = 9'h18f == r_count_56_io_out ? io_r_399_b : _GEN_22978; // @[SWChisel.scala 221:{19,19}]
  assign array_56_io_e_i = E_56; // @[SWChisel.scala 196:21]
  assign array_56_io_f_i = F_56; // @[SWChisel.scala 198:21]
  assign array_56_io_ve_i = V1_57; // @[SWChisel.scala 197:22]
  assign array_56_io_vf_i = V1_56; // @[SWChisel.scala 199:22]
  assign array_56_io_vv_i = V2_56; // @[SWChisel.scala 200:22]
  assign array_57_io_q = io_q_57_b; // @[SWChisel.scala 220:19]
  assign array_57_io_r = 9'h18f == r_count_57_io_out ? io_r_399_b : _GEN_23378; // @[SWChisel.scala 221:{19,19}]
  assign array_57_io_e_i = E_57; // @[SWChisel.scala 196:21]
  assign array_57_io_f_i = F_57; // @[SWChisel.scala 198:21]
  assign array_57_io_ve_i = V1_58; // @[SWChisel.scala 197:22]
  assign array_57_io_vf_i = V1_57; // @[SWChisel.scala 199:22]
  assign array_57_io_vv_i = V2_57; // @[SWChisel.scala 200:22]
  assign array_58_io_q = io_q_58_b; // @[SWChisel.scala 220:19]
  assign array_58_io_r = 9'h18f == r_count_58_io_out ? io_r_399_b : _GEN_23778; // @[SWChisel.scala 221:{19,19}]
  assign array_58_io_e_i = E_58; // @[SWChisel.scala 196:21]
  assign array_58_io_f_i = F_58; // @[SWChisel.scala 198:21]
  assign array_58_io_ve_i = V1_59; // @[SWChisel.scala 197:22]
  assign array_58_io_vf_i = V1_58; // @[SWChisel.scala 199:22]
  assign array_58_io_vv_i = V2_58; // @[SWChisel.scala 200:22]
  assign array_59_io_q = io_q_59_b; // @[SWChisel.scala 220:19]
  assign array_59_io_r = 9'h18f == r_count_59_io_out ? io_r_399_b : _GEN_24178; // @[SWChisel.scala 221:{19,19}]
  assign array_59_io_e_i = E_59; // @[SWChisel.scala 196:21]
  assign array_59_io_f_i = F_59; // @[SWChisel.scala 198:21]
  assign array_59_io_ve_i = V1_60; // @[SWChisel.scala 197:22]
  assign array_59_io_vf_i = V1_59; // @[SWChisel.scala 199:22]
  assign array_59_io_vv_i = V2_59; // @[SWChisel.scala 200:22]
  assign r_count_0_clock = clock;
  assign r_count_0_reset = reset;
  assign r_count_0_io_en = start_reg_0; // @[SWChisel.scala 192:22]
  assign r_count_1_clock = clock;
  assign r_count_1_reset = reset;
  assign r_count_1_io_en = start_reg_1; // @[SWChisel.scala 192:22]
  assign r_count_2_clock = clock;
  assign r_count_2_reset = reset;
  assign r_count_2_io_en = start_reg_2; // @[SWChisel.scala 192:22]
  assign r_count_3_clock = clock;
  assign r_count_3_reset = reset;
  assign r_count_3_io_en = start_reg_3; // @[SWChisel.scala 192:22]
  assign r_count_4_clock = clock;
  assign r_count_4_reset = reset;
  assign r_count_4_io_en = start_reg_4; // @[SWChisel.scala 192:22]
  assign r_count_5_clock = clock;
  assign r_count_5_reset = reset;
  assign r_count_5_io_en = start_reg_5; // @[SWChisel.scala 192:22]
  assign r_count_6_clock = clock;
  assign r_count_6_reset = reset;
  assign r_count_6_io_en = start_reg_6; // @[SWChisel.scala 192:22]
  assign r_count_7_clock = clock;
  assign r_count_7_reset = reset;
  assign r_count_7_io_en = start_reg_7; // @[SWChisel.scala 192:22]
  assign r_count_8_clock = clock;
  assign r_count_8_reset = reset;
  assign r_count_8_io_en = start_reg_8; // @[SWChisel.scala 192:22]
  assign r_count_9_clock = clock;
  assign r_count_9_reset = reset;
  assign r_count_9_io_en = start_reg_9; // @[SWChisel.scala 192:22]
  assign r_count_10_clock = clock;
  assign r_count_10_reset = reset;
  assign r_count_10_io_en = start_reg_10; // @[SWChisel.scala 192:22]
  assign r_count_11_clock = clock;
  assign r_count_11_reset = reset;
  assign r_count_11_io_en = start_reg_11; // @[SWChisel.scala 192:22]
  assign r_count_12_clock = clock;
  assign r_count_12_reset = reset;
  assign r_count_12_io_en = start_reg_12; // @[SWChisel.scala 192:22]
  assign r_count_13_clock = clock;
  assign r_count_13_reset = reset;
  assign r_count_13_io_en = start_reg_13; // @[SWChisel.scala 192:22]
  assign r_count_14_clock = clock;
  assign r_count_14_reset = reset;
  assign r_count_14_io_en = start_reg_14; // @[SWChisel.scala 192:22]
  assign r_count_15_clock = clock;
  assign r_count_15_reset = reset;
  assign r_count_15_io_en = start_reg_15; // @[SWChisel.scala 192:22]
  assign r_count_16_clock = clock;
  assign r_count_16_reset = reset;
  assign r_count_16_io_en = start_reg_16; // @[SWChisel.scala 192:22]
  assign r_count_17_clock = clock;
  assign r_count_17_reset = reset;
  assign r_count_17_io_en = start_reg_17; // @[SWChisel.scala 192:22]
  assign r_count_18_clock = clock;
  assign r_count_18_reset = reset;
  assign r_count_18_io_en = start_reg_18; // @[SWChisel.scala 192:22]
  assign r_count_19_clock = clock;
  assign r_count_19_reset = reset;
  assign r_count_19_io_en = start_reg_19; // @[SWChisel.scala 192:22]
  assign r_count_20_clock = clock;
  assign r_count_20_reset = reset;
  assign r_count_20_io_en = start_reg_20; // @[SWChisel.scala 192:22]
  assign r_count_21_clock = clock;
  assign r_count_21_reset = reset;
  assign r_count_21_io_en = start_reg_21; // @[SWChisel.scala 192:22]
  assign r_count_22_clock = clock;
  assign r_count_22_reset = reset;
  assign r_count_22_io_en = start_reg_22; // @[SWChisel.scala 192:22]
  assign r_count_23_clock = clock;
  assign r_count_23_reset = reset;
  assign r_count_23_io_en = start_reg_23; // @[SWChisel.scala 192:22]
  assign r_count_24_clock = clock;
  assign r_count_24_reset = reset;
  assign r_count_24_io_en = start_reg_24; // @[SWChisel.scala 192:22]
  assign r_count_25_clock = clock;
  assign r_count_25_reset = reset;
  assign r_count_25_io_en = start_reg_25; // @[SWChisel.scala 192:22]
  assign r_count_26_clock = clock;
  assign r_count_26_reset = reset;
  assign r_count_26_io_en = start_reg_26; // @[SWChisel.scala 192:22]
  assign r_count_27_clock = clock;
  assign r_count_27_reset = reset;
  assign r_count_27_io_en = start_reg_27; // @[SWChisel.scala 192:22]
  assign r_count_28_clock = clock;
  assign r_count_28_reset = reset;
  assign r_count_28_io_en = start_reg_28; // @[SWChisel.scala 192:22]
  assign r_count_29_clock = clock;
  assign r_count_29_reset = reset;
  assign r_count_29_io_en = start_reg_29; // @[SWChisel.scala 192:22]
  assign r_count_30_clock = clock;
  assign r_count_30_reset = reset;
  assign r_count_30_io_en = start_reg_30; // @[SWChisel.scala 192:22]
  assign r_count_31_clock = clock;
  assign r_count_31_reset = reset;
  assign r_count_31_io_en = start_reg_31; // @[SWChisel.scala 192:22]
  assign r_count_32_clock = clock;
  assign r_count_32_reset = reset;
  assign r_count_32_io_en = start_reg_32; // @[SWChisel.scala 192:22]
  assign r_count_33_clock = clock;
  assign r_count_33_reset = reset;
  assign r_count_33_io_en = start_reg_33; // @[SWChisel.scala 192:22]
  assign r_count_34_clock = clock;
  assign r_count_34_reset = reset;
  assign r_count_34_io_en = start_reg_34; // @[SWChisel.scala 192:22]
  assign r_count_35_clock = clock;
  assign r_count_35_reset = reset;
  assign r_count_35_io_en = start_reg_35; // @[SWChisel.scala 192:22]
  assign r_count_36_clock = clock;
  assign r_count_36_reset = reset;
  assign r_count_36_io_en = start_reg_36; // @[SWChisel.scala 192:22]
  assign r_count_37_clock = clock;
  assign r_count_37_reset = reset;
  assign r_count_37_io_en = start_reg_37; // @[SWChisel.scala 192:22]
  assign r_count_38_clock = clock;
  assign r_count_38_reset = reset;
  assign r_count_38_io_en = start_reg_38; // @[SWChisel.scala 192:22]
  assign r_count_39_clock = clock;
  assign r_count_39_reset = reset;
  assign r_count_39_io_en = start_reg_39; // @[SWChisel.scala 192:22]
  assign r_count_40_clock = clock;
  assign r_count_40_reset = reset;
  assign r_count_40_io_en = start_reg_40; // @[SWChisel.scala 192:22]
  assign r_count_41_clock = clock;
  assign r_count_41_reset = reset;
  assign r_count_41_io_en = start_reg_41; // @[SWChisel.scala 192:22]
  assign r_count_42_clock = clock;
  assign r_count_42_reset = reset;
  assign r_count_42_io_en = start_reg_42; // @[SWChisel.scala 192:22]
  assign r_count_43_clock = clock;
  assign r_count_43_reset = reset;
  assign r_count_43_io_en = start_reg_43; // @[SWChisel.scala 192:22]
  assign r_count_44_clock = clock;
  assign r_count_44_reset = reset;
  assign r_count_44_io_en = start_reg_44; // @[SWChisel.scala 192:22]
  assign r_count_45_clock = clock;
  assign r_count_45_reset = reset;
  assign r_count_45_io_en = start_reg_45; // @[SWChisel.scala 192:22]
  assign r_count_46_clock = clock;
  assign r_count_46_reset = reset;
  assign r_count_46_io_en = start_reg_46; // @[SWChisel.scala 192:22]
  assign r_count_47_clock = clock;
  assign r_count_47_reset = reset;
  assign r_count_47_io_en = start_reg_47; // @[SWChisel.scala 192:22]
  assign r_count_48_clock = clock;
  assign r_count_48_reset = reset;
  assign r_count_48_io_en = start_reg_48; // @[SWChisel.scala 192:22]
  assign r_count_49_clock = clock;
  assign r_count_49_reset = reset;
  assign r_count_49_io_en = start_reg_49; // @[SWChisel.scala 192:22]
  assign r_count_50_clock = clock;
  assign r_count_50_reset = reset;
  assign r_count_50_io_en = start_reg_50; // @[SWChisel.scala 192:22]
  assign r_count_51_clock = clock;
  assign r_count_51_reset = reset;
  assign r_count_51_io_en = start_reg_51; // @[SWChisel.scala 192:22]
  assign r_count_52_clock = clock;
  assign r_count_52_reset = reset;
  assign r_count_52_io_en = start_reg_52; // @[SWChisel.scala 192:22]
  assign r_count_53_clock = clock;
  assign r_count_53_reset = reset;
  assign r_count_53_io_en = start_reg_53; // @[SWChisel.scala 192:22]
  assign r_count_54_clock = clock;
  assign r_count_54_reset = reset;
  assign r_count_54_io_en = start_reg_54; // @[SWChisel.scala 192:22]
  assign r_count_55_clock = clock;
  assign r_count_55_reset = reset;
  assign r_count_55_io_en = start_reg_55; // @[SWChisel.scala 192:22]
  assign r_count_56_clock = clock;
  assign r_count_56_reset = reset;
  assign r_count_56_io_en = start_reg_56; // @[SWChisel.scala 192:22]
  assign r_count_57_clock = clock;
  assign r_count_57_reset = reset;
  assign r_count_57_io_en = start_reg_57; // @[SWChisel.scala 192:22]
  assign r_count_58_clock = clock;
  assign r_count_58_reset = reset;
  assign r_count_58_io_en = start_reg_58; // @[SWChisel.scala 192:22]
  assign r_count_59_clock = clock;
  assign r_count_59_reset = reset;
  assign r_count_59_io_en = start_reg_59; // @[SWChisel.scala 192:22]
  assign max_clock = clock;
  assign max_reset = reset;
  assign max_io_start = start_reg_59; // @[SWChisel.scala 178:16]
  assign max_io_in = V1_60; // @[SWChisel.scala 177:13]
  always @(posedge clock) begin
    if (reset) begin // @[SWChisel.scala 162:18]
      E_0 <= -16'sh2; // @[SWChisel.scala 162:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      E_0 <= array_0_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_1 <= -16'sh3; // @[SWChisel.scala 162:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      E_1 <= array_1_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_2 <= -16'sh4; // @[SWChisel.scala 162:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      E_2 <= array_2_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_3 <= -16'sh5; // @[SWChisel.scala 162:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      E_3 <= array_3_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_4 <= -16'sh6; // @[SWChisel.scala 162:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      E_4 <= array_4_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_5 <= -16'sh7; // @[SWChisel.scala 162:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      E_5 <= array_5_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_6 <= -16'sh8; // @[SWChisel.scala 162:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      E_6 <= array_6_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_7 <= -16'sh9; // @[SWChisel.scala 162:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      E_7 <= array_7_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_8 <= -16'sha; // @[SWChisel.scala 162:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      E_8 <= array_8_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_9 <= -16'shb; // @[SWChisel.scala 162:18]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      E_9 <= array_9_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_10 <= -16'shc; // @[SWChisel.scala 162:18]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      E_10 <= array_10_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_11 <= -16'shd; // @[SWChisel.scala 162:18]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      E_11 <= array_11_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_12 <= -16'she; // @[SWChisel.scala 162:18]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      E_12 <= array_12_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_13 <= -16'shf; // @[SWChisel.scala 162:18]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      E_13 <= array_13_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_14 <= -16'sh10; // @[SWChisel.scala 162:18]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      E_14 <= array_14_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_15 <= -16'sh11; // @[SWChisel.scala 162:18]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      E_15 <= array_15_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_16 <= -16'sh12; // @[SWChisel.scala 162:18]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      E_16 <= array_16_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_17 <= -16'sh13; // @[SWChisel.scala 162:18]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      E_17 <= array_17_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_18 <= -16'sh14; // @[SWChisel.scala 162:18]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      E_18 <= array_18_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_19 <= -16'sh15; // @[SWChisel.scala 162:18]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      E_19 <= array_19_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_20 <= -16'sh16; // @[SWChisel.scala 162:18]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      E_20 <= array_20_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_21 <= -16'sh17; // @[SWChisel.scala 162:18]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      E_21 <= array_21_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_22 <= -16'sh18; // @[SWChisel.scala 162:18]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      E_22 <= array_22_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_23 <= -16'sh19; // @[SWChisel.scala 162:18]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      E_23 <= array_23_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_24 <= -16'sh1a; // @[SWChisel.scala 162:18]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      E_24 <= array_24_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_25 <= -16'sh1b; // @[SWChisel.scala 162:18]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      E_25 <= array_25_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_26 <= -16'sh1c; // @[SWChisel.scala 162:18]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      E_26 <= array_26_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_27 <= -16'sh1d; // @[SWChisel.scala 162:18]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      E_27 <= array_27_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_28 <= -16'sh1e; // @[SWChisel.scala 162:18]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      E_28 <= array_28_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_29 <= -16'sh1f; // @[SWChisel.scala 162:18]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      E_29 <= array_29_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_30 <= -16'sh20; // @[SWChisel.scala 162:18]
    end else if (start_reg_30) begin // @[SWChisel.scala 207:25]
      E_30 <= array_30_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_31 <= -16'sh21; // @[SWChisel.scala 162:18]
    end else if (start_reg_31) begin // @[SWChisel.scala 207:25]
      E_31 <= array_31_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_32 <= -16'sh22; // @[SWChisel.scala 162:18]
    end else if (start_reg_32) begin // @[SWChisel.scala 207:25]
      E_32 <= array_32_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_33 <= -16'sh23; // @[SWChisel.scala 162:18]
    end else if (start_reg_33) begin // @[SWChisel.scala 207:25]
      E_33 <= array_33_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_34 <= -16'sh24; // @[SWChisel.scala 162:18]
    end else if (start_reg_34) begin // @[SWChisel.scala 207:25]
      E_34 <= array_34_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_35 <= -16'sh25; // @[SWChisel.scala 162:18]
    end else if (start_reg_35) begin // @[SWChisel.scala 207:25]
      E_35 <= array_35_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_36 <= -16'sh26; // @[SWChisel.scala 162:18]
    end else if (start_reg_36) begin // @[SWChisel.scala 207:25]
      E_36 <= array_36_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_37 <= -16'sh27; // @[SWChisel.scala 162:18]
    end else if (start_reg_37) begin // @[SWChisel.scala 207:25]
      E_37 <= array_37_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_38 <= -16'sh28; // @[SWChisel.scala 162:18]
    end else if (start_reg_38) begin // @[SWChisel.scala 207:25]
      E_38 <= array_38_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_39 <= -16'sh29; // @[SWChisel.scala 162:18]
    end else if (start_reg_39) begin // @[SWChisel.scala 207:25]
      E_39 <= array_39_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_40 <= -16'sh2a; // @[SWChisel.scala 162:18]
    end else if (start_reg_40) begin // @[SWChisel.scala 207:25]
      E_40 <= array_40_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_41 <= -16'sh2b; // @[SWChisel.scala 162:18]
    end else if (start_reg_41) begin // @[SWChisel.scala 207:25]
      E_41 <= array_41_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_42 <= -16'sh2c; // @[SWChisel.scala 162:18]
    end else if (start_reg_42) begin // @[SWChisel.scala 207:25]
      E_42 <= array_42_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_43 <= -16'sh2d; // @[SWChisel.scala 162:18]
    end else if (start_reg_43) begin // @[SWChisel.scala 207:25]
      E_43 <= array_43_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_44 <= -16'sh2e; // @[SWChisel.scala 162:18]
    end else if (start_reg_44) begin // @[SWChisel.scala 207:25]
      E_44 <= array_44_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_45 <= -16'sh2f; // @[SWChisel.scala 162:18]
    end else if (start_reg_45) begin // @[SWChisel.scala 207:25]
      E_45 <= array_45_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_46 <= -16'sh30; // @[SWChisel.scala 162:18]
    end else if (start_reg_46) begin // @[SWChisel.scala 207:25]
      E_46 <= array_46_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_47 <= -16'sh31; // @[SWChisel.scala 162:18]
    end else if (start_reg_47) begin // @[SWChisel.scala 207:25]
      E_47 <= array_47_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_48 <= -16'sh32; // @[SWChisel.scala 162:18]
    end else if (start_reg_48) begin // @[SWChisel.scala 207:25]
      E_48 <= array_48_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_49 <= -16'sh33; // @[SWChisel.scala 162:18]
    end else if (start_reg_49) begin // @[SWChisel.scala 207:25]
      E_49 <= array_49_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_50 <= -16'sh34; // @[SWChisel.scala 162:18]
    end else if (start_reg_50) begin // @[SWChisel.scala 207:25]
      E_50 <= array_50_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_51 <= -16'sh35; // @[SWChisel.scala 162:18]
    end else if (start_reg_51) begin // @[SWChisel.scala 207:25]
      E_51 <= array_51_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_52 <= -16'sh36; // @[SWChisel.scala 162:18]
    end else if (start_reg_52) begin // @[SWChisel.scala 207:25]
      E_52 <= array_52_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_53 <= -16'sh37; // @[SWChisel.scala 162:18]
    end else if (start_reg_53) begin // @[SWChisel.scala 207:25]
      E_53 <= array_53_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_54 <= -16'sh38; // @[SWChisel.scala 162:18]
    end else if (start_reg_54) begin // @[SWChisel.scala 207:25]
      E_54 <= array_54_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_55 <= -16'sh39; // @[SWChisel.scala 162:18]
    end else if (start_reg_55) begin // @[SWChisel.scala 207:25]
      E_55 <= array_55_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_56 <= -16'sh3a; // @[SWChisel.scala 162:18]
    end else if (start_reg_56) begin // @[SWChisel.scala 207:25]
      E_56 <= array_56_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_57 <= -16'sh3b; // @[SWChisel.scala 162:18]
    end else if (start_reg_57) begin // @[SWChisel.scala 207:25]
      E_57 <= array_57_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_58 <= -16'sh3c; // @[SWChisel.scala 162:18]
    end else if (start_reg_58) begin // @[SWChisel.scala 207:25]
      E_58 <= array_58_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_59 <= -16'sh3d; // @[SWChisel.scala 162:18]
    end else if (start_reg_59) begin // @[SWChisel.scala 207:25]
      E_59 <= array_59_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_1 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      F_1 <= array_0_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_2 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      F_2 <= array_1_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_3 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      F_3 <= array_2_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_4 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      F_4 <= array_3_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_5 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      F_5 <= array_4_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_6 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      F_6 <= array_5_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_7 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      F_7 <= array_6_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_8 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      F_8 <= array_7_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_9 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      F_9 <= array_8_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_10 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      F_10 <= array_9_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_11 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      F_11 <= array_10_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_12 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      F_12 <= array_11_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_13 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      F_13 <= array_12_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_14 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      F_14 <= array_13_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_15 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      F_15 <= array_14_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_16 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      F_16 <= array_15_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_17 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      F_17 <= array_16_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_18 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      F_18 <= array_17_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_19 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      F_19 <= array_18_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_20 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      F_20 <= array_19_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_21 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      F_21 <= array_20_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_22 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      F_22 <= array_21_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_23 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      F_23 <= array_22_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_24 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      F_24 <= array_23_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_25 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      F_25 <= array_24_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_26 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      F_26 <= array_25_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_27 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      F_27 <= array_26_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_28 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      F_28 <= array_27_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_29 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      F_29 <= array_28_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_30 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      F_30 <= array_29_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_31 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_30) begin // @[SWChisel.scala 207:25]
      F_31 <= array_30_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_32 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_31) begin // @[SWChisel.scala 207:25]
      F_32 <= array_31_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_33 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_32) begin // @[SWChisel.scala 207:25]
      F_33 <= array_32_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_34 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_33) begin // @[SWChisel.scala 207:25]
      F_34 <= array_33_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_35 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_34) begin // @[SWChisel.scala 207:25]
      F_35 <= array_34_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_36 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_35) begin // @[SWChisel.scala 207:25]
      F_36 <= array_35_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_37 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_36) begin // @[SWChisel.scala 207:25]
      F_37 <= array_36_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_38 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_37) begin // @[SWChisel.scala 207:25]
      F_38 <= array_37_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_39 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_38) begin // @[SWChisel.scala 207:25]
      F_39 <= array_38_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_40 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_39) begin // @[SWChisel.scala 207:25]
      F_40 <= array_39_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_41 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_40) begin // @[SWChisel.scala 207:25]
      F_41 <= array_40_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_42 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_41) begin // @[SWChisel.scala 207:25]
      F_42 <= array_41_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_43 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_42) begin // @[SWChisel.scala 207:25]
      F_43 <= array_42_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_44 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_43) begin // @[SWChisel.scala 207:25]
      F_44 <= array_43_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_45 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_44) begin // @[SWChisel.scala 207:25]
      F_45 <= array_44_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_46 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_45) begin // @[SWChisel.scala 207:25]
      F_46 <= array_45_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_47 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_46) begin // @[SWChisel.scala 207:25]
      F_47 <= array_46_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_48 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_47) begin // @[SWChisel.scala 207:25]
      F_48 <= array_47_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_49 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_48) begin // @[SWChisel.scala 207:25]
      F_49 <= array_48_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_50 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_49) begin // @[SWChisel.scala 207:25]
      F_50 <= array_49_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_51 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_50) begin // @[SWChisel.scala 207:25]
      F_51 <= array_50_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_52 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_51) begin // @[SWChisel.scala 207:25]
      F_52 <= array_51_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_53 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_52) begin // @[SWChisel.scala 207:25]
      F_53 <= array_52_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_54 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_53) begin // @[SWChisel.scala 207:25]
      F_54 <= array_53_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_55 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_54) begin // @[SWChisel.scala 207:25]
      F_55 <= array_54_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_56 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_55) begin // @[SWChisel.scala 207:25]
      F_56 <= array_55_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_57 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_56) begin // @[SWChisel.scala 207:25]
      F_57 <= array_56_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_58 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_57) begin // @[SWChisel.scala 207:25]
      F_58 <= array_57_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_59 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_58) begin // @[SWChisel.scala 207:25]
      F_59 <= array_58_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_0 <= -16'sh1; // @[SWChisel.scala 164:19]
    end else begin
      V1_0 <= 16'sh0; // @[SWChisel.scala 165:9]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_1 <= -16'sh2; // @[SWChisel.scala 164:19]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      V1_1 <= array_0_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_2 <= -16'sh3; // @[SWChisel.scala 164:19]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      V1_2 <= array_1_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_3 <= -16'sh4; // @[SWChisel.scala 164:19]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      V1_3 <= array_2_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_4 <= -16'sh5; // @[SWChisel.scala 164:19]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      V1_4 <= array_3_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_5 <= -16'sh6; // @[SWChisel.scala 164:19]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      V1_5 <= array_4_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_6 <= -16'sh7; // @[SWChisel.scala 164:19]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      V1_6 <= array_5_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_7 <= -16'sh8; // @[SWChisel.scala 164:19]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      V1_7 <= array_6_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_8 <= -16'sh9; // @[SWChisel.scala 164:19]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      V1_8 <= array_7_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_9 <= -16'sha; // @[SWChisel.scala 164:19]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      V1_9 <= array_8_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_10 <= -16'shb; // @[SWChisel.scala 164:19]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      V1_10 <= array_9_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_11 <= -16'shc; // @[SWChisel.scala 164:19]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      V1_11 <= array_10_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_12 <= -16'shd; // @[SWChisel.scala 164:19]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      V1_12 <= array_11_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_13 <= -16'she; // @[SWChisel.scala 164:19]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      V1_13 <= array_12_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_14 <= -16'shf; // @[SWChisel.scala 164:19]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      V1_14 <= array_13_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_15 <= -16'sh10; // @[SWChisel.scala 164:19]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      V1_15 <= array_14_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_16 <= -16'sh11; // @[SWChisel.scala 164:19]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      V1_16 <= array_15_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_17 <= -16'sh12; // @[SWChisel.scala 164:19]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      V1_17 <= array_16_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_18 <= -16'sh13; // @[SWChisel.scala 164:19]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      V1_18 <= array_17_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_19 <= -16'sh14; // @[SWChisel.scala 164:19]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      V1_19 <= array_18_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_20 <= -16'sh15; // @[SWChisel.scala 164:19]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      V1_20 <= array_19_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_21 <= -16'sh16; // @[SWChisel.scala 164:19]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      V1_21 <= array_20_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_22 <= -16'sh17; // @[SWChisel.scala 164:19]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      V1_22 <= array_21_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_23 <= -16'sh18; // @[SWChisel.scala 164:19]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      V1_23 <= array_22_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_24 <= -16'sh19; // @[SWChisel.scala 164:19]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      V1_24 <= array_23_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_25 <= -16'sh1a; // @[SWChisel.scala 164:19]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      V1_25 <= array_24_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_26 <= -16'sh1b; // @[SWChisel.scala 164:19]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      V1_26 <= array_25_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_27 <= -16'sh1c; // @[SWChisel.scala 164:19]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      V1_27 <= array_26_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_28 <= -16'sh1d; // @[SWChisel.scala 164:19]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      V1_28 <= array_27_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_29 <= -16'sh1e; // @[SWChisel.scala 164:19]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      V1_29 <= array_28_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_30 <= -16'sh1f; // @[SWChisel.scala 164:19]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      V1_30 <= array_29_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_31 <= -16'sh20; // @[SWChisel.scala 164:19]
    end else if (start_reg_30) begin // @[SWChisel.scala 207:25]
      V1_31 <= array_30_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_32 <= -16'sh21; // @[SWChisel.scala 164:19]
    end else if (start_reg_31) begin // @[SWChisel.scala 207:25]
      V1_32 <= array_31_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_33 <= -16'sh22; // @[SWChisel.scala 164:19]
    end else if (start_reg_32) begin // @[SWChisel.scala 207:25]
      V1_33 <= array_32_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_34 <= -16'sh23; // @[SWChisel.scala 164:19]
    end else if (start_reg_33) begin // @[SWChisel.scala 207:25]
      V1_34 <= array_33_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_35 <= -16'sh24; // @[SWChisel.scala 164:19]
    end else if (start_reg_34) begin // @[SWChisel.scala 207:25]
      V1_35 <= array_34_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_36 <= -16'sh25; // @[SWChisel.scala 164:19]
    end else if (start_reg_35) begin // @[SWChisel.scala 207:25]
      V1_36 <= array_35_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_37 <= -16'sh26; // @[SWChisel.scala 164:19]
    end else if (start_reg_36) begin // @[SWChisel.scala 207:25]
      V1_37 <= array_36_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_38 <= -16'sh27; // @[SWChisel.scala 164:19]
    end else if (start_reg_37) begin // @[SWChisel.scala 207:25]
      V1_38 <= array_37_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_39 <= -16'sh28; // @[SWChisel.scala 164:19]
    end else if (start_reg_38) begin // @[SWChisel.scala 207:25]
      V1_39 <= array_38_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_40 <= -16'sh29; // @[SWChisel.scala 164:19]
    end else if (start_reg_39) begin // @[SWChisel.scala 207:25]
      V1_40 <= array_39_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_41 <= -16'sh2a; // @[SWChisel.scala 164:19]
    end else if (start_reg_40) begin // @[SWChisel.scala 207:25]
      V1_41 <= array_40_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_42 <= -16'sh2b; // @[SWChisel.scala 164:19]
    end else if (start_reg_41) begin // @[SWChisel.scala 207:25]
      V1_42 <= array_41_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_43 <= -16'sh2c; // @[SWChisel.scala 164:19]
    end else if (start_reg_42) begin // @[SWChisel.scala 207:25]
      V1_43 <= array_42_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_44 <= -16'sh2d; // @[SWChisel.scala 164:19]
    end else if (start_reg_43) begin // @[SWChisel.scala 207:25]
      V1_44 <= array_43_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_45 <= -16'sh2e; // @[SWChisel.scala 164:19]
    end else if (start_reg_44) begin // @[SWChisel.scala 207:25]
      V1_45 <= array_44_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_46 <= -16'sh2f; // @[SWChisel.scala 164:19]
    end else if (start_reg_45) begin // @[SWChisel.scala 207:25]
      V1_46 <= array_45_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_47 <= -16'sh30; // @[SWChisel.scala 164:19]
    end else if (start_reg_46) begin // @[SWChisel.scala 207:25]
      V1_47 <= array_46_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_48 <= -16'sh31; // @[SWChisel.scala 164:19]
    end else if (start_reg_47) begin // @[SWChisel.scala 207:25]
      V1_48 <= array_47_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_49 <= -16'sh32; // @[SWChisel.scala 164:19]
    end else if (start_reg_48) begin // @[SWChisel.scala 207:25]
      V1_49 <= array_48_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_50 <= -16'sh33; // @[SWChisel.scala 164:19]
    end else if (start_reg_49) begin // @[SWChisel.scala 207:25]
      V1_50 <= array_49_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_51 <= -16'sh34; // @[SWChisel.scala 164:19]
    end else if (start_reg_50) begin // @[SWChisel.scala 207:25]
      V1_51 <= array_50_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_52 <= -16'sh35; // @[SWChisel.scala 164:19]
    end else if (start_reg_51) begin // @[SWChisel.scala 207:25]
      V1_52 <= array_51_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_53 <= -16'sh36; // @[SWChisel.scala 164:19]
    end else if (start_reg_52) begin // @[SWChisel.scala 207:25]
      V1_53 <= array_52_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_54 <= -16'sh37; // @[SWChisel.scala 164:19]
    end else if (start_reg_53) begin // @[SWChisel.scala 207:25]
      V1_54 <= array_53_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_55 <= -16'sh38; // @[SWChisel.scala 164:19]
    end else if (start_reg_54) begin // @[SWChisel.scala 207:25]
      V1_55 <= array_54_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_56 <= -16'sh39; // @[SWChisel.scala 164:19]
    end else if (start_reg_55) begin // @[SWChisel.scala 207:25]
      V1_56 <= array_55_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_57 <= -16'sh3a; // @[SWChisel.scala 164:19]
    end else if (start_reg_56) begin // @[SWChisel.scala 207:25]
      V1_57 <= array_56_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_58 <= -16'sh3b; // @[SWChisel.scala 164:19]
    end else if (start_reg_57) begin // @[SWChisel.scala 207:25]
      V1_58 <= array_57_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_59 <= -16'sh3c; // @[SWChisel.scala 164:19]
    end else if (start_reg_58) begin // @[SWChisel.scala 207:25]
      V1_59 <= array_58_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_60 <= -16'sh3d; // @[SWChisel.scala 164:19]
    end else if (start_reg_59) begin // @[SWChisel.scala 207:25]
      V1_60 <= array_59_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_0 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_0 <= V1_0; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_1 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_1 <= V1_1; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_2 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_2 <= V1_2; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_3 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_3 <= V1_3; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_4 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_4 <= V1_4; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_5 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_5 <= V1_5; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_6 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_6 <= V1_6; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_7 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_7 <= V1_7; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_8 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_8 <= V1_8; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_9 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_9 <= V1_9; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_10 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_10 <= V1_10; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_11 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_11 <= V1_11; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_12 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_12 <= V1_12; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_13 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_13 <= V1_13; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_14 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_14 <= V1_14; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_15 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_15 <= V1_15; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_16 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_16 <= V1_16; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_17 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_17 <= V1_17; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_18 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_18 <= V1_18; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_19 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_19 <= V1_19; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_20 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_20 <= V1_20; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_21 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_21 <= V1_21; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_22 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_22 <= V1_22; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_23 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_23 <= V1_23; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_24 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_24 <= V1_24; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_25 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_25 <= V1_25; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_26 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_26 <= V1_26; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_27 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_27 <= V1_27; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_28 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_28 <= V1_28; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_29 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_29 <= V1_29; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_30 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_30 <= V1_30; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_31 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_31 <= V1_31; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_32 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_32 <= V1_32; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_33 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_33 <= V1_33; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_34 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_34 <= V1_34; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_35 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_35 <= V1_35; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_36 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_36 <= V1_36; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_37 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_37 <= V1_37; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_38 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_38 <= V1_38; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_39 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_39 <= V1_39; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_40 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_40 <= V1_40; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_41 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_41 <= V1_41; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_42 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_42 <= V1_42; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_43 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_43 <= V1_43; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_44 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_44 <= V1_44; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_45 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_45 <= V1_45; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_46 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_46 <= V1_46; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_47 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_47 <= V1_47; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_48 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_48 <= V1_48; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_49 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_49 <= V1_49; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_50 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_50 <= V1_50; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_51 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_51 <= V1_51; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_52 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_52 <= V1_52; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_53 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_53 <= V1_53; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_54 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_54 <= V1_54; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_55 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_55 <= V1_55; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_56 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_56 <= V1_56; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_57 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_57 <= V1_57; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_58 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_58 <= V1_58; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_59 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_59 <= V1_59; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_0 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_0 <= io_start; // @[SWChisel.scala 185:16]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_1 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_1 <= start_reg_0; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_2 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_2 <= start_reg_1; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_3 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_3 <= start_reg_2; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_4 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_4 <= start_reg_3; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_5 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_5 <= start_reg_4; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_6 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_6 <= start_reg_5; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_7 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_7 <= start_reg_6; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_8 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_8 <= start_reg_7; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_9 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_9 <= start_reg_8; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_10 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_10 <= start_reg_9; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_11 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_11 <= start_reg_10; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_12 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_12 <= start_reg_11; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_13 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_13 <= start_reg_12; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_14 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_14 <= start_reg_13; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_15 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_15 <= start_reg_14; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_16 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_16 <= start_reg_15; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_17 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_17 <= start_reg_16; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_18 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_18 <= start_reg_17; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_19 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_19 <= start_reg_18; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_20 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_20 <= start_reg_19; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_21 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_21 <= start_reg_20; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_22 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_22 <= start_reg_21; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_23 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_23 <= start_reg_22; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_24 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_24 <= start_reg_23; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_25 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_25 <= start_reg_24; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_26 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_26 <= start_reg_25; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_27 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_27 <= start_reg_26; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_28 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_28 <= start_reg_27; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_29 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_29 <= start_reg_28; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_30 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_30 <= start_reg_29; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_31 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_31 <= start_reg_30; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_32 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_32 <= start_reg_31; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_33 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_33 <= start_reg_32; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_34 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_34 <= start_reg_33; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_35 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_35 <= start_reg_34; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_36 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_36 <= start_reg_35; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_37 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_37 <= start_reg_36; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_38 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_38 <= start_reg_37; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_39 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_39 <= start_reg_38; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_40 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_40 <= start_reg_39; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_41 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_41 <= start_reg_40; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_42 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_42 <= start_reg_41; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_43 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_43 <= start_reg_42; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_44 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_44 <= start_reg_43; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_45 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_45 <= start_reg_44; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_46 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_46 <= start_reg_45; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_47 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_47 <= start_reg_46; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_48 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_48 <= start_reg_47; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_49 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_49 <= start_reg_48; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_50 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_50 <= start_reg_49; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_51 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_51 <= start_reg_50; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_52 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_52 <= start_reg_51; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_53 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_53 <= start_reg_52; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_54 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_54 <= start_reg_53; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_55 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_55 <= start_reg_54; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_56 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_56 <= start_reg_55; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_57 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_57 <= start_reg_56; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_58 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_58 <= start_reg_57; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_59 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_59 <= start_reg_58; // @[SWChisel.scala 187:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  E_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  E_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  E_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  E_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  E_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  E_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  E_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  E_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  E_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  E_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  E_10 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  E_11 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  E_12 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  E_13 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  E_14 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  E_15 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  E_16 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  E_17 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  E_18 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  E_19 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  E_20 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  E_21 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  E_22 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  E_23 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  E_24 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  E_25 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  E_26 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  E_27 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  E_28 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  E_29 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  E_30 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  E_31 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  E_32 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  E_33 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  E_34 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  E_35 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  E_36 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  E_37 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  E_38 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  E_39 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  E_40 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  E_41 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  E_42 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  E_43 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  E_44 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  E_45 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  E_46 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  E_47 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  E_48 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  E_49 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  E_50 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  E_51 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  E_52 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  E_53 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  E_54 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  E_55 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  E_56 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  E_57 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  E_58 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  E_59 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  F_1 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  F_2 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  F_3 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  F_4 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  F_5 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  F_6 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  F_7 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  F_8 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  F_9 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  F_10 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  F_11 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  F_12 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  F_13 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  F_14 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  F_15 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  F_16 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  F_17 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  F_18 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  F_19 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  F_20 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  F_21 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  F_22 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  F_23 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  F_24 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  F_25 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  F_26 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  F_27 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  F_28 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  F_29 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  F_30 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  F_31 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  F_32 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  F_33 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  F_34 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  F_35 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  F_36 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  F_37 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  F_38 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  F_39 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  F_40 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  F_41 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  F_42 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  F_43 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  F_44 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  F_45 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  F_46 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  F_47 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  F_48 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  F_49 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  F_50 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  F_51 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  F_52 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  F_53 = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  F_54 = _RAND_113[15:0];
  _RAND_114 = {1{`RANDOM}};
  F_55 = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  F_56 = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  F_57 = _RAND_116[15:0];
  _RAND_117 = {1{`RANDOM}};
  F_58 = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  F_59 = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  V1_0 = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  V1_1 = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  V1_2 = _RAND_121[15:0];
  _RAND_122 = {1{`RANDOM}};
  V1_3 = _RAND_122[15:0];
  _RAND_123 = {1{`RANDOM}};
  V1_4 = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  V1_5 = _RAND_124[15:0];
  _RAND_125 = {1{`RANDOM}};
  V1_6 = _RAND_125[15:0];
  _RAND_126 = {1{`RANDOM}};
  V1_7 = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  V1_8 = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  V1_9 = _RAND_128[15:0];
  _RAND_129 = {1{`RANDOM}};
  V1_10 = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  V1_11 = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  V1_12 = _RAND_131[15:0];
  _RAND_132 = {1{`RANDOM}};
  V1_13 = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  V1_14 = _RAND_133[15:0];
  _RAND_134 = {1{`RANDOM}};
  V1_15 = _RAND_134[15:0];
  _RAND_135 = {1{`RANDOM}};
  V1_16 = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  V1_17 = _RAND_136[15:0];
  _RAND_137 = {1{`RANDOM}};
  V1_18 = _RAND_137[15:0];
  _RAND_138 = {1{`RANDOM}};
  V1_19 = _RAND_138[15:0];
  _RAND_139 = {1{`RANDOM}};
  V1_20 = _RAND_139[15:0];
  _RAND_140 = {1{`RANDOM}};
  V1_21 = _RAND_140[15:0];
  _RAND_141 = {1{`RANDOM}};
  V1_22 = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  V1_23 = _RAND_142[15:0];
  _RAND_143 = {1{`RANDOM}};
  V1_24 = _RAND_143[15:0];
  _RAND_144 = {1{`RANDOM}};
  V1_25 = _RAND_144[15:0];
  _RAND_145 = {1{`RANDOM}};
  V1_26 = _RAND_145[15:0];
  _RAND_146 = {1{`RANDOM}};
  V1_27 = _RAND_146[15:0];
  _RAND_147 = {1{`RANDOM}};
  V1_28 = _RAND_147[15:0];
  _RAND_148 = {1{`RANDOM}};
  V1_29 = _RAND_148[15:0];
  _RAND_149 = {1{`RANDOM}};
  V1_30 = _RAND_149[15:0];
  _RAND_150 = {1{`RANDOM}};
  V1_31 = _RAND_150[15:0];
  _RAND_151 = {1{`RANDOM}};
  V1_32 = _RAND_151[15:0];
  _RAND_152 = {1{`RANDOM}};
  V1_33 = _RAND_152[15:0];
  _RAND_153 = {1{`RANDOM}};
  V1_34 = _RAND_153[15:0];
  _RAND_154 = {1{`RANDOM}};
  V1_35 = _RAND_154[15:0];
  _RAND_155 = {1{`RANDOM}};
  V1_36 = _RAND_155[15:0];
  _RAND_156 = {1{`RANDOM}};
  V1_37 = _RAND_156[15:0];
  _RAND_157 = {1{`RANDOM}};
  V1_38 = _RAND_157[15:0];
  _RAND_158 = {1{`RANDOM}};
  V1_39 = _RAND_158[15:0];
  _RAND_159 = {1{`RANDOM}};
  V1_40 = _RAND_159[15:0];
  _RAND_160 = {1{`RANDOM}};
  V1_41 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  V1_42 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  V1_43 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  V1_44 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  V1_45 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  V1_46 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  V1_47 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  V1_48 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  V1_49 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  V1_50 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  V1_51 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  V1_52 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  V1_53 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  V1_54 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  V1_55 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  V1_56 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  V1_57 = _RAND_176[15:0];
  _RAND_177 = {1{`RANDOM}};
  V1_58 = _RAND_177[15:0];
  _RAND_178 = {1{`RANDOM}};
  V1_59 = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  V1_60 = _RAND_179[15:0];
  _RAND_180 = {1{`RANDOM}};
  V2_0 = _RAND_180[15:0];
  _RAND_181 = {1{`RANDOM}};
  V2_1 = _RAND_181[15:0];
  _RAND_182 = {1{`RANDOM}};
  V2_2 = _RAND_182[15:0];
  _RAND_183 = {1{`RANDOM}};
  V2_3 = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  V2_4 = _RAND_184[15:0];
  _RAND_185 = {1{`RANDOM}};
  V2_5 = _RAND_185[15:0];
  _RAND_186 = {1{`RANDOM}};
  V2_6 = _RAND_186[15:0];
  _RAND_187 = {1{`RANDOM}};
  V2_7 = _RAND_187[15:0];
  _RAND_188 = {1{`RANDOM}};
  V2_8 = _RAND_188[15:0];
  _RAND_189 = {1{`RANDOM}};
  V2_9 = _RAND_189[15:0];
  _RAND_190 = {1{`RANDOM}};
  V2_10 = _RAND_190[15:0];
  _RAND_191 = {1{`RANDOM}};
  V2_11 = _RAND_191[15:0];
  _RAND_192 = {1{`RANDOM}};
  V2_12 = _RAND_192[15:0];
  _RAND_193 = {1{`RANDOM}};
  V2_13 = _RAND_193[15:0];
  _RAND_194 = {1{`RANDOM}};
  V2_14 = _RAND_194[15:0];
  _RAND_195 = {1{`RANDOM}};
  V2_15 = _RAND_195[15:0];
  _RAND_196 = {1{`RANDOM}};
  V2_16 = _RAND_196[15:0];
  _RAND_197 = {1{`RANDOM}};
  V2_17 = _RAND_197[15:0];
  _RAND_198 = {1{`RANDOM}};
  V2_18 = _RAND_198[15:0];
  _RAND_199 = {1{`RANDOM}};
  V2_19 = _RAND_199[15:0];
  _RAND_200 = {1{`RANDOM}};
  V2_20 = _RAND_200[15:0];
  _RAND_201 = {1{`RANDOM}};
  V2_21 = _RAND_201[15:0];
  _RAND_202 = {1{`RANDOM}};
  V2_22 = _RAND_202[15:0];
  _RAND_203 = {1{`RANDOM}};
  V2_23 = _RAND_203[15:0];
  _RAND_204 = {1{`RANDOM}};
  V2_24 = _RAND_204[15:0];
  _RAND_205 = {1{`RANDOM}};
  V2_25 = _RAND_205[15:0];
  _RAND_206 = {1{`RANDOM}};
  V2_26 = _RAND_206[15:0];
  _RAND_207 = {1{`RANDOM}};
  V2_27 = _RAND_207[15:0];
  _RAND_208 = {1{`RANDOM}};
  V2_28 = _RAND_208[15:0];
  _RAND_209 = {1{`RANDOM}};
  V2_29 = _RAND_209[15:0];
  _RAND_210 = {1{`RANDOM}};
  V2_30 = _RAND_210[15:0];
  _RAND_211 = {1{`RANDOM}};
  V2_31 = _RAND_211[15:0];
  _RAND_212 = {1{`RANDOM}};
  V2_32 = _RAND_212[15:0];
  _RAND_213 = {1{`RANDOM}};
  V2_33 = _RAND_213[15:0];
  _RAND_214 = {1{`RANDOM}};
  V2_34 = _RAND_214[15:0];
  _RAND_215 = {1{`RANDOM}};
  V2_35 = _RAND_215[15:0];
  _RAND_216 = {1{`RANDOM}};
  V2_36 = _RAND_216[15:0];
  _RAND_217 = {1{`RANDOM}};
  V2_37 = _RAND_217[15:0];
  _RAND_218 = {1{`RANDOM}};
  V2_38 = _RAND_218[15:0];
  _RAND_219 = {1{`RANDOM}};
  V2_39 = _RAND_219[15:0];
  _RAND_220 = {1{`RANDOM}};
  V2_40 = _RAND_220[15:0];
  _RAND_221 = {1{`RANDOM}};
  V2_41 = _RAND_221[15:0];
  _RAND_222 = {1{`RANDOM}};
  V2_42 = _RAND_222[15:0];
  _RAND_223 = {1{`RANDOM}};
  V2_43 = _RAND_223[15:0];
  _RAND_224 = {1{`RANDOM}};
  V2_44 = _RAND_224[15:0];
  _RAND_225 = {1{`RANDOM}};
  V2_45 = _RAND_225[15:0];
  _RAND_226 = {1{`RANDOM}};
  V2_46 = _RAND_226[15:0];
  _RAND_227 = {1{`RANDOM}};
  V2_47 = _RAND_227[15:0];
  _RAND_228 = {1{`RANDOM}};
  V2_48 = _RAND_228[15:0];
  _RAND_229 = {1{`RANDOM}};
  V2_49 = _RAND_229[15:0];
  _RAND_230 = {1{`RANDOM}};
  V2_50 = _RAND_230[15:0];
  _RAND_231 = {1{`RANDOM}};
  V2_51 = _RAND_231[15:0];
  _RAND_232 = {1{`RANDOM}};
  V2_52 = _RAND_232[15:0];
  _RAND_233 = {1{`RANDOM}};
  V2_53 = _RAND_233[15:0];
  _RAND_234 = {1{`RANDOM}};
  V2_54 = _RAND_234[15:0];
  _RAND_235 = {1{`RANDOM}};
  V2_55 = _RAND_235[15:0];
  _RAND_236 = {1{`RANDOM}};
  V2_56 = _RAND_236[15:0];
  _RAND_237 = {1{`RANDOM}};
  V2_57 = _RAND_237[15:0];
  _RAND_238 = {1{`RANDOM}};
  V2_58 = _RAND_238[15:0];
  _RAND_239 = {1{`RANDOM}};
  V2_59 = _RAND_239[15:0];
  _RAND_240 = {1{`RANDOM}};
  start_reg_0 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  start_reg_1 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  start_reg_2 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  start_reg_3 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  start_reg_4 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  start_reg_5 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  start_reg_6 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  start_reg_7 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  start_reg_8 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  start_reg_9 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  start_reg_10 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  start_reg_11 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  start_reg_12 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  start_reg_13 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  start_reg_14 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  start_reg_15 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  start_reg_16 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  start_reg_17 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  start_reg_18 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  start_reg_19 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  start_reg_20 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  start_reg_21 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  start_reg_22 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  start_reg_23 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  start_reg_24 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  start_reg_25 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  start_reg_26 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  start_reg_27 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  start_reg_28 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  start_reg_29 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  start_reg_30 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  start_reg_31 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  start_reg_32 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  start_reg_33 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  start_reg_34 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  start_reg_35 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  start_reg_36 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  start_reg_37 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  start_reg_38 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  start_reg_39 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  start_reg_40 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  start_reg_41 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  start_reg_42 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  start_reg_43 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  start_reg_44 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  start_reg_45 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  start_reg_46 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  start_reg_47 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  start_reg_48 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  start_reg_49 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  start_reg_50 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  start_reg_51 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  start_reg_52 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  start_reg_53 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  start_reg_54 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  start_reg_55 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  start_reg_56 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  start_reg_57 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  start_reg_58 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  start_reg_59 = _RAND_299[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
