module SWCell(
  input  [1:0]  io_q,
  input  [1:0]  io_r,
  input  [15:0] io_e_i,
  input  [15:0] io_f_i,
  input  [15:0] io_ve_i,
  input  [15:0] io_vf_i,
  input  [15:0] io_vv_i,
  output [15:0] io_e_o,
  output [15:0] io_f_o,
  output [15:0] io_v_o
);
  wire [15:0] _T_2 = $signed(io_ve_i) - 16'sh2; // @[SWChisel.scala 78:17]
  wire [15:0] _T_5 = $signed(io_e_i) - 16'sh1; // @[SWChisel.scala 78:39]
  wire [15:0] e_max = $signed(_T_2) >= $signed(_T_5) ? $signed(_T_2) : $signed(_T_5); // @[SWChisel.scala 78:51 79:11 81:11]
  wire [15:0] _T_9 = $signed(io_vf_i) - 16'sh2; // @[SWChisel.scala 85:17]
  wire [15:0] _T_12 = $signed(io_f_i) - 16'sh1; // @[SWChisel.scala 85:38]
  wire [15:0] f_max = $signed(_T_9) > $signed(_T_12) ? $signed(_T_9) : $signed(_T_12); // @[SWChisel.scala 85:50 86:11 88:11]
  wire [15:0] ef_temp = $signed(e_max) > $signed(f_max) ? $signed(e_max) : $signed(f_max); // @[SWChisel.scala 92:24 93:13 95:13]
  wire [15:0] _v_temp_T_2 = $signed(io_vv_i) + 16'sh2; // @[SWChisel.scala 100:23]
  wire [15:0] _v_temp_T_5 = $signed(io_vv_i) - 16'sh2; // @[SWChisel.scala 102:23]
  wire [15:0] v_temp = io_q == io_r ? $signed(_v_temp_T_2) : $signed(_v_temp_T_5); // @[SWChisel.scala 100:12 102:12 99:24]
  assign io_e_o = $signed(_T_2) >= $signed(_T_5) ? $signed(_T_2) : $signed(_T_5); // @[SWChisel.scala 78:51 79:11 81:11]
  assign io_f_o = $signed(_T_9) > $signed(_T_12) ? $signed(_T_9) : $signed(_T_12); // @[SWChisel.scala 85:50 86:11 88:11]
  assign io_v_o = $signed(v_temp) > $signed(ef_temp) ? $signed(v_temp) : $signed(ef_temp); // @[SWChisel.scala 106:27 107:11 109:11]
endmodule
module MyCounter(
  input        clock,
  input        reset,
  input        io_en,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [6:0] _io_out_T_2 = io_out + 7'h1; // @[SWChisel.scala 155:55]
  reg [6:0] io_out_r; // @[Reg.scala 35:20]
  assign io_out = io_out_r; // @[SWChisel.scala 155:12]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      io_out_r <= 7'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_out < 7'h64) begin // @[SWChisel.scala 155:28]
        io_out_r <= _io_out_T_2;
      end else begin
        io_out_r <= 7'h0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_out_r = _RAND_0[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MAX(
  input         clock,
  input         reset,
  input         io_start,
  input  [15:0] io_in,
  output        io_done,
  output [15:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] max; // @[SWChisel.scala 122:20]
  reg [6:0] counter; // @[SWChisel.scala 133:24]
  wire [6:0] _counter_T_1 = counter - 7'h1; // @[SWChisel.scala 135:24]
  assign io_done = counter == 7'h0; // @[SWChisel.scala 141:17]
  assign io_out = max; // @[SWChisel.scala 123:10]
  always @(posedge clock) begin
    if (reset) begin // @[SWChisel.scala 122:20]
      max <= 16'sh8000; // @[SWChisel.scala 122:20]
    end else if ($signed(io_in) > $signed(max)) begin // @[SWChisel.scala 126:22]
      max <= io_in; // @[SWChisel.scala 127:9]
    end
    if (reset) begin // @[SWChisel.scala 133:24]
      counter <= 7'h65; // @[SWChisel.scala 133:24]
    end else if (counter == 7'h0) begin // @[SWChisel.scala 141:26]
      counter <= 7'h0; // @[SWChisel.scala 143:13]
    end else if (io_start) begin // @[SWChisel.scala 134:19]
      counter <= _counter_T_1; // @[SWChisel.scala 135:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  max = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SW(
  input         clock,
  input         reset,
  input  [1:0]  io_q_0_b,
  input  [1:0]  io_q_1_b,
  input  [1:0]  io_q_2_b,
  input  [1:0]  io_q_3_b,
  input  [1:0]  io_q_4_b,
  input  [1:0]  io_q_5_b,
  input  [1:0]  io_q_6_b,
  input  [1:0]  io_q_7_b,
  input  [1:0]  io_q_8_b,
  input  [1:0]  io_q_9_b,
  input  [1:0]  io_r_0_b,
  input  [1:0]  io_r_1_b,
  input  [1:0]  io_r_2_b,
  input  [1:0]  io_r_3_b,
  input  [1:0]  io_r_4_b,
  input  [1:0]  io_r_5_b,
  input  [1:0]  io_r_6_b,
  input  [1:0]  io_r_7_b,
  input  [1:0]  io_r_8_b,
  input  [1:0]  io_r_9_b,
  input  [1:0]  io_r_10_b,
  input  [1:0]  io_r_11_b,
  input  [1:0]  io_r_12_b,
  input  [1:0]  io_r_13_b,
  input  [1:0]  io_r_14_b,
  input  [1:0]  io_r_15_b,
  input  [1:0]  io_r_16_b,
  input  [1:0]  io_r_17_b,
  input  [1:0]  io_r_18_b,
  input  [1:0]  io_r_19_b,
  input  [1:0]  io_r_20_b,
  input  [1:0]  io_r_21_b,
  input  [1:0]  io_r_22_b,
  input  [1:0]  io_r_23_b,
  input  [1:0]  io_r_24_b,
  input  [1:0]  io_r_25_b,
  input  [1:0]  io_r_26_b,
  input  [1:0]  io_r_27_b,
  input  [1:0]  io_r_28_b,
  input  [1:0]  io_r_29_b,
  input  [1:0]  io_r_30_b,
  input  [1:0]  io_r_31_b,
  input  [1:0]  io_r_32_b,
  input  [1:0]  io_r_33_b,
  input  [1:0]  io_r_34_b,
  input  [1:0]  io_r_35_b,
  input  [1:0]  io_r_36_b,
  input  [1:0]  io_r_37_b,
  input  [1:0]  io_r_38_b,
  input  [1:0]  io_r_39_b,
  input  [1:0]  io_r_40_b,
  input  [1:0]  io_r_41_b,
  input  [1:0]  io_r_42_b,
  input  [1:0]  io_r_43_b,
  input  [1:0]  io_r_44_b,
  input  [1:0]  io_r_45_b,
  input  [1:0]  io_r_46_b,
  input  [1:0]  io_r_47_b,
  input  [1:0]  io_r_48_b,
  input  [1:0]  io_r_49_b,
  input  [1:0]  io_r_50_b,
  input  [1:0]  io_r_51_b,
  input  [1:0]  io_r_52_b,
  input  [1:0]  io_r_53_b,
  input  [1:0]  io_r_54_b,
  input  [1:0]  io_r_55_b,
  input  [1:0]  io_r_56_b,
  input  [1:0]  io_r_57_b,
  input  [1:0]  io_r_58_b,
  input  [1:0]  io_r_59_b,
  input  [1:0]  io_r_60_b,
  input  [1:0]  io_r_61_b,
  input  [1:0]  io_r_62_b,
  input  [1:0]  io_r_63_b,
  input  [1:0]  io_r_64_b,
  input  [1:0]  io_r_65_b,
  input  [1:0]  io_r_66_b,
  input  [1:0]  io_r_67_b,
  input  [1:0]  io_r_68_b,
  input  [1:0]  io_r_69_b,
  input  [1:0]  io_r_70_b,
  input  [1:0]  io_r_71_b,
  input  [1:0]  io_r_72_b,
  input  [1:0]  io_r_73_b,
  input  [1:0]  io_r_74_b,
  input  [1:0]  io_r_75_b,
  input  [1:0]  io_r_76_b,
  input  [1:0]  io_r_77_b,
  input  [1:0]  io_r_78_b,
  input  [1:0]  io_r_79_b,
  input  [1:0]  io_r_80_b,
  input  [1:0]  io_r_81_b,
  input  [1:0]  io_r_82_b,
  input  [1:0]  io_r_83_b,
  input  [1:0]  io_r_84_b,
  input  [1:0]  io_r_85_b,
  input  [1:0]  io_r_86_b,
  input  [1:0]  io_r_87_b,
  input  [1:0]  io_r_88_b,
  input  [1:0]  io_r_89_b,
  input  [1:0]  io_r_90_b,
  input  [1:0]  io_r_91_b,
  input  [1:0]  io_r_92_b,
  input  [1:0]  io_r_93_b,
  input  [1:0]  io_r_94_b,
  input  [1:0]  io_r_95_b,
  input  [1:0]  io_r_96_b,
  input  [1:0]  io_r_97_b,
  input  [1:0]  io_r_98_b,
  input  [1:0]  io_r_99_b,
  input         io_start,
  output [15:0] io_result,
  output        io_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] array_0_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_0_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_1_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_1_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_2_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_2_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_3_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_3_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_4_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_4_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_5_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_5_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_6_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_6_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_7_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_7_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_8_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_8_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_9_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_9_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_v_o; // @[SWChisel.scala 170:39]
  wire  r_count_0_clock; // @[SWChisel.scala 171:41]
  wire  r_count_0_reset; // @[SWChisel.scala 171:41]
  wire  r_count_0_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_0_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_1_clock; // @[SWChisel.scala 171:41]
  wire  r_count_1_reset; // @[SWChisel.scala 171:41]
  wire  r_count_1_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_1_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_2_clock; // @[SWChisel.scala 171:41]
  wire  r_count_2_reset; // @[SWChisel.scala 171:41]
  wire  r_count_2_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_2_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_3_clock; // @[SWChisel.scala 171:41]
  wire  r_count_3_reset; // @[SWChisel.scala 171:41]
  wire  r_count_3_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_3_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_4_clock; // @[SWChisel.scala 171:41]
  wire  r_count_4_reset; // @[SWChisel.scala 171:41]
  wire  r_count_4_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_4_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_5_clock; // @[SWChisel.scala 171:41]
  wire  r_count_5_reset; // @[SWChisel.scala 171:41]
  wire  r_count_5_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_5_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_6_clock; // @[SWChisel.scala 171:41]
  wire  r_count_6_reset; // @[SWChisel.scala 171:41]
  wire  r_count_6_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_6_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_7_clock; // @[SWChisel.scala 171:41]
  wire  r_count_7_reset; // @[SWChisel.scala 171:41]
  wire  r_count_7_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_7_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_8_clock; // @[SWChisel.scala 171:41]
  wire  r_count_8_reset; // @[SWChisel.scala 171:41]
  wire  r_count_8_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_8_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_9_clock; // @[SWChisel.scala 171:41]
  wire  r_count_9_reset; // @[SWChisel.scala 171:41]
  wire  r_count_9_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_9_io_out; // @[SWChisel.scala 171:41]
  wire  max_clock; // @[SWChisel.scala 174:19]
  wire  max_reset; // @[SWChisel.scala 174:19]
  wire  max_io_start; // @[SWChisel.scala 174:19]
  wire [15:0] max_io_in; // @[SWChisel.scala 174:19]
  wire  max_io_done; // @[SWChisel.scala 174:19]
  wire [15:0] max_io_out; // @[SWChisel.scala 174:19]
  reg [15:0] E_0; // @[SWChisel.scala 162:18]
  reg [15:0] E_1; // @[SWChisel.scala 162:18]
  reg [15:0] E_2; // @[SWChisel.scala 162:18]
  reg [15:0] E_3; // @[SWChisel.scala 162:18]
  reg [15:0] E_4; // @[SWChisel.scala 162:18]
  reg [15:0] E_5; // @[SWChisel.scala 162:18]
  reg [15:0] E_6; // @[SWChisel.scala 162:18]
  reg [15:0] E_7; // @[SWChisel.scala 162:18]
  reg [15:0] E_8; // @[SWChisel.scala 162:18]
  reg [15:0] E_9; // @[SWChisel.scala 162:18]
  reg [15:0] F_1; // @[SWChisel.scala 163:18]
  reg [15:0] F_2; // @[SWChisel.scala 163:18]
  reg [15:0] F_3; // @[SWChisel.scala 163:18]
  reg [15:0] F_4; // @[SWChisel.scala 163:18]
  reg [15:0] F_5; // @[SWChisel.scala 163:18]
  reg [15:0] F_6; // @[SWChisel.scala 163:18]
  reg [15:0] F_7; // @[SWChisel.scala 163:18]
  reg [15:0] F_8; // @[SWChisel.scala 163:18]
  reg [15:0] F_9; // @[SWChisel.scala 163:18]
  reg [15:0] V1_0; // @[SWChisel.scala 164:19]
  reg [15:0] V1_1; // @[SWChisel.scala 164:19]
  reg [15:0] V1_2; // @[SWChisel.scala 164:19]
  reg [15:0] V1_3; // @[SWChisel.scala 164:19]
  reg [15:0] V1_4; // @[SWChisel.scala 164:19]
  reg [15:0] V1_5; // @[SWChisel.scala 164:19]
  reg [15:0] V1_6; // @[SWChisel.scala 164:19]
  reg [15:0] V1_7; // @[SWChisel.scala 164:19]
  reg [15:0] V1_8; // @[SWChisel.scala 164:19]
  reg [15:0] V1_9; // @[SWChisel.scala 164:19]
  reg [15:0] V1_10; // @[SWChisel.scala 164:19]
  reg [15:0] V2_0; // @[SWChisel.scala 166:19]
  reg [15:0] V2_1; // @[SWChisel.scala 166:19]
  reg [15:0] V2_2; // @[SWChisel.scala 166:19]
  reg [15:0] V2_3; // @[SWChisel.scala 166:19]
  reg [15:0] V2_4; // @[SWChisel.scala 166:19]
  reg [15:0] V2_5; // @[SWChisel.scala 166:19]
  reg [15:0] V2_6; // @[SWChisel.scala 166:19]
  reg [15:0] V2_7; // @[SWChisel.scala 166:19]
  reg [15:0] V2_8; // @[SWChisel.scala 166:19]
  reg [15:0] V2_9; // @[SWChisel.scala 166:19]
  reg  start_reg_0; // @[SWChisel.scala 167:26]
  reg  start_reg_1; // @[SWChisel.scala 167:26]
  reg  start_reg_2; // @[SWChisel.scala 167:26]
  reg  start_reg_3; // @[SWChisel.scala 167:26]
  reg  start_reg_4; // @[SWChisel.scala 167:26]
  reg  start_reg_5; // @[SWChisel.scala 167:26]
  reg  start_reg_6; // @[SWChisel.scala 167:26]
  reg  start_reg_7; // @[SWChisel.scala 167:26]
  reg  start_reg_8; // @[SWChisel.scala 167:26]
  reg  start_reg_9; // @[SWChisel.scala 167:26]
  wire [1:0] _GEN_31 = 7'h1 == r_count_0_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_32 = 7'h2 == r_count_0_io_out ? io_r_2_b : _GEN_31; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_33 = 7'h3 == r_count_0_io_out ? io_r_3_b : _GEN_32; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_34 = 7'h4 == r_count_0_io_out ? io_r_4_b : _GEN_33; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_35 = 7'h5 == r_count_0_io_out ? io_r_5_b : _GEN_34; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_36 = 7'h6 == r_count_0_io_out ? io_r_6_b : _GEN_35; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_37 = 7'h7 == r_count_0_io_out ? io_r_7_b : _GEN_36; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_38 = 7'h8 == r_count_0_io_out ? io_r_8_b : _GEN_37; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_39 = 7'h9 == r_count_0_io_out ? io_r_9_b : _GEN_38; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_40 = 7'ha == r_count_0_io_out ? io_r_10_b : _GEN_39; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_41 = 7'hb == r_count_0_io_out ? io_r_11_b : _GEN_40; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_42 = 7'hc == r_count_0_io_out ? io_r_12_b : _GEN_41; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_43 = 7'hd == r_count_0_io_out ? io_r_13_b : _GEN_42; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_44 = 7'he == r_count_0_io_out ? io_r_14_b : _GEN_43; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_45 = 7'hf == r_count_0_io_out ? io_r_15_b : _GEN_44; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_46 = 7'h10 == r_count_0_io_out ? io_r_16_b : _GEN_45; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_47 = 7'h11 == r_count_0_io_out ? io_r_17_b : _GEN_46; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_48 = 7'h12 == r_count_0_io_out ? io_r_18_b : _GEN_47; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_49 = 7'h13 == r_count_0_io_out ? io_r_19_b : _GEN_48; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_50 = 7'h14 == r_count_0_io_out ? io_r_20_b : _GEN_49; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_51 = 7'h15 == r_count_0_io_out ? io_r_21_b : _GEN_50; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_52 = 7'h16 == r_count_0_io_out ? io_r_22_b : _GEN_51; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_53 = 7'h17 == r_count_0_io_out ? io_r_23_b : _GEN_52; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_54 = 7'h18 == r_count_0_io_out ? io_r_24_b : _GEN_53; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_55 = 7'h19 == r_count_0_io_out ? io_r_25_b : _GEN_54; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_56 = 7'h1a == r_count_0_io_out ? io_r_26_b : _GEN_55; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_57 = 7'h1b == r_count_0_io_out ? io_r_27_b : _GEN_56; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_58 = 7'h1c == r_count_0_io_out ? io_r_28_b : _GEN_57; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_59 = 7'h1d == r_count_0_io_out ? io_r_29_b : _GEN_58; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_60 = 7'h1e == r_count_0_io_out ? io_r_30_b : _GEN_59; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_61 = 7'h1f == r_count_0_io_out ? io_r_31_b : _GEN_60; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_62 = 7'h20 == r_count_0_io_out ? io_r_32_b : _GEN_61; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_63 = 7'h21 == r_count_0_io_out ? io_r_33_b : _GEN_62; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_64 = 7'h22 == r_count_0_io_out ? io_r_34_b : _GEN_63; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_65 = 7'h23 == r_count_0_io_out ? io_r_35_b : _GEN_64; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_66 = 7'h24 == r_count_0_io_out ? io_r_36_b : _GEN_65; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_67 = 7'h25 == r_count_0_io_out ? io_r_37_b : _GEN_66; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_68 = 7'h26 == r_count_0_io_out ? io_r_38_b : _GEN_67; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_69 = 7'h27 == r_count_0_io_out ? io_r_39_b : _GEN_68; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_70 = 7'h28 == r_count_0_io_out ? io_r_40_b : _GEN_69; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_71 = 7'h29 == r_count_0_io_out ? io_r_41_b : _GEN_70; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_72 = 7'h2a == r_count_0_io_out ? io_r_42_b : _GEN_71; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_73 = 7'h2b == r_count_0_io_out ? io_r_43_b : _GEN_72; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_74 = 7'h2c == r_count_0_io_out ? io_r_44_b : _GEN_73; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_75 = 7'h2d == r_count_0_io_out ? io_r_45_b : _GEN_74; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_76 = 7'h2e == r_count_0_io_out ? io_r_46_b : _GEN_75; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_77 = 7'h2f == r_count_0_io_out ? io_r_47_b : _GEN_76; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_78 = 7'h30 == r_count_0_io_out ? io_r_48_b : _GEN_77; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_79 = 7'h31 == r_count_0_io_out ? io_r_49_b : _GEN_78; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_80 = 7'h32 == r_count_0_io_out ? io_r_50_b : _GEN_79; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_81 = 7'h33 == r_count_0_io_out ? io_r_51_b : _GEN_80; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_82 = 7'h34 == r_count_0_io_out ? io_r_52_b : _GEN_81; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_83 = 7'h35 == r_count_0_io_out ? io_r_53_b : _GEN_82; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_84 = 7'h36 == r_count_0_io_out ? io_r_54_b : _GEN_83; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_85 = 7'h37 == r_count_0_io_out ? io_r_55_b : _GEN_84; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_86 = 7'h38 == r_count_0_io_out ? io_r_56_b : _GEN_85; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_87 = 7'h39 == r_count_0_io_out ? io_r_57_b : _GEN_86; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_88 = 7'h3a == r_count_0_io_out ? io_r_58_b : _GEN_87; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_89 = 7'h3b == r_count_0_io_out ? io_r_59_b : _GEN_88; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_90 = 7'h3c == r_count_0_io_out ? io_r_60_b : _GEN_89; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_91 = 7'h3d == r_count_0_io_out ? io_r_61_b : _GEN_90; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_92 = 7'h3e == r_count_0_io_out ? io_r_62_b : _GEN_91; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_93 = 7'h3f == r_count_0_io_out ? io_r_63_b : _GEN_92; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_94 = 7'h40 == r_count_0_io_out ? io_r_64_b : _GEN_93; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_95 = 7'h41 == r_count_0_io_out ? io_r_65_b : _GEN_94; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_96 = 7'h42 == r_count_0_io_out ? io_r_66_b : _GEN_95; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_97 = 7'h43 == r_count_0_io_out ? io_r_67_b : _GEN_96; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_98 = 7'h44 == r_count_0_io_out ? io_r_68_b : _GEN_97; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_99 = 7'h45 == r_count_0_io_out ? io_r_69_b : _GEN_98; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_100 = 7'h46 == r_count_0_io_out ? io_r_70_b : _GEN_99; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_101 = 7'h47 == r_count_0_io_out ? io_r_71_b : _GEN_100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_102 = 7'h48 == r_count_0_io_out ? io_r_72_b : _GEN_101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_103 = 7'h49 == r_count_0_io_out ? io_r_73_b : _GEN_102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_104 = 7'h4a == r_count_0_io_out ? io_r_74_b : _GEN_103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_105 = 7'h4b == r_count_0_io_out ? io_r_75_b : _GEN_104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_106 = 7'h4c == r_count_0_io_out ? io_r_76_b : _GEN_105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_107 = 7'h4d == r_count_0_io_out ? io_r_77_b : _GEN_106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_108 = 7'h4e == r_count_0_io_out ? io_r_78_b : _GEN_107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_109 = 7'h4f == r_count_0_io_out ? io_r_79_b : _GEN_108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_110 = 7'h50 == r_count_0_io_out ? io_r_80_b : _GEN_109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_111 = 7'h51 == r_count_0_io_out ? io_r_81_b : _GEN_110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_112 = 7'h52 == r_count_0_io_out ? io_r_82_b : _GEN_111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_113 = 7'h53 == r_count_0_io_out ? io_r_83_b : _GEN_112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_114 = 7'h54 == r_count_0_io_out ? io_r_84_b : _GEN_113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_115 = 7'h55 == r_count_0_io_out ? io_r_85_b : _GEN_114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_116 = 7'h56 == r_count_0_io_out ? io_r_86_b : _GEN_115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_117 = 7'h57 == r_count_0_io_out ? io_r_87_b : _GEN_116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_118 = 7'h58 == r_count_0_io_out ? io_r_88_b : _GEN_117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_119 = 7'h59 == r_count_0_io_out ? io_r_89_b : _GEN_118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_120 = 7'h5a == r_count_0_io_out ? io_r_90_b : _GEN_119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_121 = 7'h5b == r_count_0_io_out ? io_r_91_b : _GEN_120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_122 = 7'h5c == r_count_0_io_out ? io_r_92_b : _GEN_121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_123 = 7'h5d == r_count_0_io_out ? io_r_93_b : _GEN_122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_124 = 7'h5e == r_count_0_io_out ? io_r_94_b : _GEN_123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_125 = 7'h5f == r_count_0_io_out ? io_r_95_b : _GEN_124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_126 = 7'h60 == r_count_0_io_out ? io_r_96_b : _GEN_125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_127 = 7'h61 == r_count_0_io_out ? io_r_97_b : _GEN_126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_128 = 7'h62 == r_count_0_io_out ? io_r_98_b : _GEN_127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_131 = 7'h1 == r_count_1_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_132 = 7'h2 == r_count_1_io_out ? io_r_2_b : _GEN_131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_133 = 7'h3 == r_count_1_io_out ? io_r_3_b : _GEN_132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_134 = 7'h4 == r_count_1_io_out ? io_r_4_b : _GEN_133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_135 = 7'h5 == r_count_1_io_out ? io_r_5_b : _GEN_134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_136 = 7'h6 == r_count_1_io_out ? io_r_6_b : _GEN_135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_137 = 7'h7 == r_count_1_io_out ? io_r_7_b : _GEN_136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_138 = 7'h8 == r_count_1_io_out ? io_r_8_b : _GEN_137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_139 = 7'h9 == r_count_1_io_out ? io_r_9_b : _GEN_138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_140 = 7'ha == r_count_1_io_out ? io_r_10_b : _GEN_139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_141 = 7'hb == r_count_1_io_out ? io_r_11_b : _GEN_140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_142 = 7'hc == r_count_1_io_out ? io_r_12_b : _GEN_141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_143 = 7'hd == r_count_1_io_out ? io_r_13_b : _GEN_142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_144 = 7'he == r_count_1_io_out ? io_r_14_b : _GEN_143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_145 = 7'hf == r_count_1_io_out ? io_r_15_b : _GEN_144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_146 = 7'h10 == r_count_1_io_out ? io_r_16_b : _GEN_145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_147 = 7'h11 == r_count_1_io_out ? io_r_17_b : _GEN_146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_148 = 7'h12 == r_count_1_io_out ? io_r_18_b : _GEN_147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_149 = 7'h13 == r_count_1_io_out ? io_r_19_b : _GEN_148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_150 = 7'h14 == r_count_1_io_out ? io_r_20_b : _GEN_149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_151 = 7'h15 == r_count_1_io_out ? io_r_21_b : _GEN_150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_152 = 7'h16 == r_count_1_io_out ? io_r_22_b : _GEN_151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_153 = 7'h17 == r_count_1_io_out ? io_r_23_b : _GEN_152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_154 = 7'h18 == r_count_1_io_out ? io_r_24_b : _GEN_153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_155 = 7'h19 == r_count_1_io_out ? io_r_25_b : _GEN_154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_156 = 7'h1a == r_count_1_io_out ? io_r_26_b : _GEN_155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_157 = 7'h1b == r_count_1_io_out ? io_r_27_b : _GEN_156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_158 = 7'h1c == r_count_1_io_out ? io_r_28_b : _GEN_157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_159 = 7'h1d == r_count_1_io_out ? io_r_29_b : _GEN_158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_160 = 7'h1e == r_count_1_io_out ? io_r_30_b : _GEN_159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_161 = 7'h1f == r_count_1_io_out ? io_r_31_b : _GEN_160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_162 = 7'h20 == r_count_1_io_out ? io_r_32_b : _GEN_161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_163 = 7'h21 == r_count_1_io_out ? io_r_33_b : _GEN_162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_164 = 7'h22 == r_count_1_io_out ? io_r_34_b : _GEN_163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_165 = 7'h23 == r_count_1_io_out ? io_r_35_b : _GEN_164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_166 = 7'h24 == r_count_1_io_out ? io_r_36_b : _GEN_165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_167 = 7'h25 == r_count_1_io_out ? io_r_37_b : _GEN_166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_168 = 7'h26 == r_count_1_io_out ? io_r_38_b : _GEN_167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_169 = 7'h27 == r_count_1_io_out ? io_r_39_b : _GEN_168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_170 = 7'h28 == r_count_1_io_out ? io_r_40_b : _GEN_169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_171 = 7'h29 == r_count_1_io_out ? io_r_41_b : _GEN_170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_172 = 7'h2a == r_count_1_io_out ? io_r_42_b : _GEN_171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_173 = 7'h2b == r_count_1_io_out ? io_r_43_b : _GEN_172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_174 = 7'h2c == r_count_1_io_out ? io_r_44_b : _GEN_173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_175 = 7'h2d == r_count_1_io_out ? io_r_45_b : _GEN_174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_176 = 7'h2e == r_count_1_io_out ? io_r_46_b : _GEN_175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_177 = 7'h2f == r_count_1_io_out ? io_r_47_b : _GEN_176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_178 = 7'h30 == r_count_1_io_out ? io_r_48_b : _GEN_177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_179 = 7'h31 == r_count_1_io_out ? io_r_49_b : _GEN_178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_180 = 7'h32 == r_count_1_io_out ? io_r_50_b : _GEN_179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_181 = 7'h33 == r_count_1_io_out ? io_r_51_b : _GEN_180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_182 = 7'h34 == r_count_1_io_out ? io_r_52_b : _GEN_181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_183 = 7'h35 == r_count_1_io_out ? io_r_53_b : _GEN_182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_184 = 7'h36 == r_count_1_io_out ? io_r_54_b : _GEN_183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_185 = 7'h37 == r_count_1_io_out ? io_r_55_b : _GEN_184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_186 = 7'h38 == r_count_1_io_out ? io_r_56_b : _GEN_185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_187 = 7'h39 == r_count_1_io_out ? io_r_57_b : _GEN_186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_188 = 7'h3a == r_count_1_io_out ? io_r_58_b : _GEN_187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_189 = 7'h3b == r_count_1_io_out ? io_r_59_b : _GEN_188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_190 = 7'h3c == r_count_1_io_out ? io_r_60_b : _GEN_189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_191 = 7'h3d == r_count_1_io_out ? io_r_61_b : _GEN_190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_192 = 7'h3e == r_count_1_io_out ? io_r_62_b : _GEN_191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_193 = 7'h3f == r_count_1_io_out ? io_r_63_b : _GEN_192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_194 = 7'h40 == r_count_1_io_out ? io_r_64_b : _GEN_193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_195 = 7'h41 == r_count_1_io_out ? io_r_65_b : _GEN_194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_196 = 7'h42 == r_count_1_io_out ? io_r_66_b : _GEN_195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_197 = 7'h43 == r_count_1_io_out ? io_r_67_b : _GEN_196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_198 = 7'h44 == r_count_1_io_out ? io_r_68_b : _GEN_197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_199 = 7'h45 == r_count_1_io_out ? io_r_69_b : _GEN_198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_200 = 7'h46 == r_count_1_io_out ? io_r_70_b : _GEN_199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_201 = 7'h47 == r_count_1_io_out ? io_r_71_b : _GEN_200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_202 = 7'h48 == r_count_1_io_out ? io_r_72_b : _GEN_201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_203 = 7'h49 == r_count_1_io_out ? io_r_73_b : _GEN_202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_204 = 7'h4a == r_count_1_io_out ? io_r_74_b : _GEN_203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_205 = 7'h4b == r_count_1_io_out ? io_r_75_b : _GEN_204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_206 = 7'h4c == r_count_1_io_out ? io_r_76_b : _GEN_205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_207 = 7'h4d == r_count_1_io_out ? io_r_77_b : _GEN_206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_208 = 7'h4e == r_count_1_io_out ? io_r_78_b : _GEN_207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_209 = 7'h4f == r_count_1_io_out ? io_r_79_b : _GEN_208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_210 = 7'h50 == r_count_1_io_out ? io_r_80_b : _GEN_209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_211 = 7'h51 == r_count_1_io_out ? io_r_81_b : _GEN_210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_212 = 7'h52 == r_count_1_io_out ? io_r_82_b : _GEN_211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_213 = 7'h53 == r_count_1_io_out ? io_r_83_b : _GEN_212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_214 = 7'h54 == r_count_1_io_out ? io_r_84_b : _GEN_213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_215 = 7'h55 == r_count_1_io_out ? io_r_85_b : _GEN_214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_216 = 7'h56 == r_count_1_io_out ? io_r_86_b : _GEN_215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_217 = 7'h57 == r_count_1_io_out ? io_r_87_b : _GEN_216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_218 = 7'h58 == r_count_1_io_out ? io_r_88_b : _GEN_217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_219 = 7'h59 == r_count_1_io_out ? io_r_89_b : _GEN_218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_220 = 7'h5a == r_count_1_io_out ? io_r_90_b : _GEN_219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_221 = 7'h5b == r_count_1_io_out ? io_r_91_b : _GEN_220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_222 = 7'h5c == r_count_1_io_out ? io_r_92_b : _GEN_221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_223 = 7'h5d == r_count_1_io_out ? io_r_93_b : _GEN_222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_224 = 7'h5e == r_count_1_io_out ? io_r_94_b : _GEN_223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_225 = 7'h5f == r_count_1_io_out ? io_r_95_b : _GEN_224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_226 = 7'h60 == r_count_1_io_out ? io_r_96_b : _GEN_225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_227 = 7'h61 == r_count_1_io_out ? io_r_97_b : _GEN_226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_228 = 7'h62 == r_count_1_io_out ? io_r_98_b : _GEN_227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_231 = 7'h1 == r_count_2_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_232 = 7'h2 == r_count_2_io_out ? io_r_2_b : _GEN_231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_233 = 7'h3 == r_count_2_io_out ? io_r_3_b : _GEN_232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_234 = 7'h4 == r_count_2_io_out ? io_r_4_b : _GEN_233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_235 = 7'h5 == r_count_2_io_out ? io_r_5_b : _GEN_234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_236 = 7'h6 == r_count_2_io_out ? io_r_6_b : _GEN_235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_237 = 7'h7 == r_count_2_io_out ? io_r_7_b : _GEN_236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_238 = 7'h8 == r_count_2_io_out ? io_r_8_b : _GEN_237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_239 = 7'h9 == r_count_2_io_out ? io_r_9_b : _GEN_238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_240 = 7'ha == r_count_2_io_out ? io_r_10_b : _GEN_239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_241 = 7'hb == r_count_2_io_out ? io_r_11_b : _GEN_240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_242 = 7'hc == r_count_2_io_out ? io_r_12_b : _GEN_241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_243 = 7'hd == r_count_2_io_out ? io_r_13_b : _GEN_242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_244 = 7'he == r_count_2_io_out ? io_r_14_b : _GEN_243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_245 = 7'hf == r_count_2_io_out ? io_r_15_b : _GEN_244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_246 = 7'h10 == r_count_2_io_out ? io_r_16_b : _GEN_245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_247 = 7'h11 == r_count_2_io_out ? io_r_17_b : _GEN_246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_248 = 7'h12 == r_count_2_io_out ? io_r_18_b : _GEN_247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_249 = 7'h13 == r_count_2_io_out ? io_r_19_b : _GEN_248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_250 = 7'h14 == r_count_2_io_out ? io_r_20_b : _GEN_249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_251 = 7'h15 == r_count_2_io_out ? io_r_21_b : _GEN_250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_252 = 7'h16 == r_count_2_io_out ? io_r_22_b : _GEN_251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_253 = 7'h17 == r_count_2_io_out ? io_r_23_b : _GEN_252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_254 = 7'h18 == r_count_2_io_out ? io_r_24_b : _GEN_253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_255 = 7'h19 == r_count_2_io_out ? io_r_25_b : _GEN_254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_256 = 7'h1a == r_count_2_io_out ? io_r_26_b : _GEN_255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_257 = 7'h1b == r_count_2_io_out ? io_r_27_b : _GEN_256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_258 = 7'h1c == r_count_2_io_out ? io_r_28_b : _GEN_257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_259 = 7'h1d == r_count_2_io_out ? io_r_29_b : _GEN_258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_260 = 7'h1e == r_count_2_io_out ? io_r_30_b : _GEN_259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_261 = 7'h1f == r_count_2_io_out ? io_r_31_b : _GEN_260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_262 = 7'h20 == r_count_2_io_out ? io_r_32_b : _GEN_261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_263 = 7'h21 == r_count_2_io_out ? io_r_33_b : _GEN_262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_264 = 7'h22 == r_count_2_io_out ? io_r_34_b : _GEN_263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_265 = 7'h23 == r_count_2_io_out ? io_r_35_b : _GEN_264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_266 = 7'h24 == r_count_2_io_out ? io_r_36_b : _GEN_265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_267 = 7'h25 == r_count_2_io_out ? io_r_37_b : _GEN_266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_268 = 7'h26 == r_count_2_io_out ? io_r_38_b : _GEN_267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_269 = 7'h27 == r_count_2_io_out ? io_r_39_b : _GEN_268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_270 = 7'h28 == r_count_2_io_out ? io_r_40_b : _GEN_269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_271 = 7'h29 == r_count_2_io_out ? io_r_41_b : _GEN_270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_272 = 7'h2a == r_count_2_io_out ? io_r_42_b : _GEN_271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_273 = 7'h2b == r_count_2_io_out ? io_r_43_b : _GEN_272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_274 = 7'h2c == r_count_2_io_out ? io_r_44_b : _GEN_273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_275 = 7'h2d == r_count_2_io_out ? io_r_45_b : _GEN_274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_276 = 7'h2e == r_count_2_io_out ? io_r_46_b : _GEN_275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_277 = 7'h2f == r_count_2_io_out ? io_r_47_b : _GEN_276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_278 = 7'h30 == r_count_2_io_out ? io_r_48_b : _GEN_277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_279 = 7'h31 == r_count_2_io_out ? io_r_49_b : _GEN_278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_280 = 7'h32 == r_count_2_io_out ? io_r_50_b : _GEN_279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_281 = 7'h33 == r_count_2_io_out ? io_r_51_b : _GEN_280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_282 = 7'h34 == r_count_2_io_out ? io_r_52_b : _GEN_281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_283 = 7'h35 == r_count_2_io_out ? io_r_53_b : _GEN_282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_284 = 7'h36 == r_count_2_io_out ? io_r_54_b : _GEN_283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_285 = 7'h37 == r_count_2_io_out ? io_r_55_b : _GEN_284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_286 = 7'h38 == r_count_2_io_out ? io_r_56_b : _GEN_285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_287 = 7'h39 == r_count_2_io_out ? io_r_57_b : _GEN_286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_288 = 7'h3a == r_count_2_io_out ? io_r_58_b : _GEN_287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_289 = 7'h3b == r_count_2_io_out ? io_r_59_b : _GEN_288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_290 = 7'h3c == r_count_2_io_out ? io_r_60_b : _GEN_289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_291 = 7'h3d == r_count_2_io_out ? io_r_61_b : _GEN_290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_292 = 7'h3e == r_count_2_io_out ? io_r_62_b : _GEN_291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_293 = 7'h3f == r_count_2_io_out ? io_r_63_b : _GEN_292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_294 = 7'h40 == r_count_2_io_out ? io_r_64_b : _GEN_293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_295 = 7'h41 == r_count_2_io_out ? io_r_65_b : _GEN_294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_296 = 7'h42 == r_count_2_io_out ? io_r_66_b : _GEN_295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_297 = 7'h43 == r_count_2_io_out ? io_r_67_b : _GEN_296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_298 = 7'h44 == r_count_2_io_out ? io_r_68_b : _GEN_297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_299 = 7'h45 == r_count_2_io_out ? io_r_69_b : _GEN_298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_300 = 7'h46 == r_count_2_io_out ? io_r_70_b : _GEN_299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_301 = 7'h47 == r_count_2_io_out ? io_r_71_b : _GEN_300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_302 = 7'h48 == r_count_2_io_out ? io_r_72_b : _GEN_301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_303 = 7'h49 == r_count_2_io_out ? io_r_73_b : _GEN_302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_304 = 7'h4a == r_count_2_io_out ? io_r_74_b : _GEN_303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_305 = 7'h4b == r_count_2_io_out ? io_r_75_b : _GEN_304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_306 = 7'h4c == r_count_2_io_out ? io_r_76_b : _GEN_305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_307 = 7'h4d == r_count_2_io_out ? io_r_77_b : _GEN_306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_308 = 7'h4e == r_count_2_io_out ? io_r_78_b : _GEN_307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_309 = 7'h4f == r_count_2_io_out ? io_r_79_b : _GEN_308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_310 = 7'h50 == r_count_2_io_out ? io_r_80_b : _GEN_309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_311 = 7'h51 == r_count_2_io_out ? io_r_81_b : _GEN_310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_312 = 7'h52 == r_count_2_io_out ? io_r_82_b : _GEN_311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_313 = 7'h53 == r_count_2_io_out ? io_r_83_b : _GEN_312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_314 = 7'h54 == r_count_2_io_out ? io_r_84_b : _GEN_313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_315 = 7'h55 == r_count_2_io_out ? io_r_85_b : _GEN_314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_316 = 7'h56 == r_count_2_io_out ? io_r_86_b : _GEN_315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_317 = 7'h57 == r_count_2_io_out ? io_r_87_b : _GEN_316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_318 = 7'h58 == r_count_2_io_out ? io_r_88_b : _GEN_317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_319 = 7'h59 == r_count_2_io_out ? io_r_89_b : _GEN_318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_320 = 7'h5a == r_count_2_io_out ? io_r_90_b : _GEN_319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_321 = 7'h5b == r_count_2_io_out ? io_r_91_b : _GEN_320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_322 = 7'h5c == r_count_2_io_out ? io_r_92_b : _GEN_321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_323 = 7'h5d == r_count_2_io_out ? io_r_93_b : _GEN_322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_324 = 7'h5e == r_count_2_io_out ? io_r_94_b : _GEN_323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_325 = 7'h5f == r_count_2_io_out ? io_r_95_b : _GEN_324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_326 = 7'h60 == r_count_2_io_out ? io_r_96_b : _GEN_325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_327 = 7'h61 == r_count_2_io_out ? io_r_97_b : _GEN_326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_328 = 7'h62 == r_count_2_io_out ? io_r_98_b : _GEN_327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_331 = 7'h1 == r_count_3_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_332 = 7'h2 == r_count_3_io_out ? io_r_2_b : _GEN_331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_333 = 7'h3 == r_count_3_io_out ? io_r_3_b : _GEN_332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_334 = 7'h4 == r_count_3_io_out ? io_r_4_b : _GEN_333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_335 = 7'h5 == r_count_3_io_out ? io_r_5_b : _GEN_334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_336 = 7'h6 == r_count_3_io_out ? io_r_6_b : _GEN_335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_337 = 7'h7 == r_count_3_io_out ? io_r_7_b : _GEN_336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_338 = 7'h8 == r_count_3_io_out ? io_r_8_b : _GEN_337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_339 = 7'h9 == r_count_3_io_out ? io_r_9_b : _GEN_338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_340 = 7'ha == r_count_3_io_out ? io_r_10_b : _GEN_339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_341 = 7'hb == r_count_3_io_out ? io_r_11_b : _GEN_340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_342 = 7'hc == r_count_3_io_out ? io_r_12_b : _GEN_341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_343 = 7'hd == r_count_3_io_out ? io_r_13_b : _GEN_342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_344 = 7'he == r_count_3_io_out ? io_r_14_b : _GEN_343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_345 = 7'hf == r_count_3_io_out ? io_r_15_b : _GEN_344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_346 = 7'h10 == r_count_3_io_out ? io_r_16_b : _GEN_345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_347 = 7'h11 == r_count_3_io_out ? io_r_17_b : _GEN_346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_348 = 7'h12 == r_count_3_io_out ? io_r_18_b : _GEN_347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_349 = 7'h13 == r_count_3_io_out ? io_r_19_b : _GEN_348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_350 = 7'h14 == r_count_3_io_out ? io_r_20_b : _GEN_349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_351 = 7'h15 == r_count_3_io_out ? io_r_21_b : _GEN_350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_352 = 7'h16 == r_count_3_io_out ? io_r_22_b : _GEN_351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_353 = 7'h17 == r_count_3_io_out ? io_r_23_b : _GEN_352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_354 = 7'h18 == r_count_3_io_out ? io_r_24_b : _GEN_353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_355 = 7'h19 == r_count_3_io_out ? io_r_25_b : _GEN_354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_356 = 7'h1a == r_count_3_io_out ? io_r_26_b : _GEN_355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_357 = 7'h1b == r_count_3_io_out ? io_r_27_b : _GEN_356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_358 = 7'h1c == r_count_3_io_out ? io_r_28_b : _GEN_357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_359 = 7'h1d == r_count_3_io_out ? io_r_29_b : _GEN_358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_360 = 7'h1e == r_count_3_io_out ? io_r_30_b : _GEN_359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_361 = 7'h1f == r_count_3_io_out ? io_r_31_b : _GEN_360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_362 = 7'h20 == r_count_3_io_out ? io_r_32_b : _GEN_361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_363 = 7'h21 == r_count_3_io_out ? io_r_33_b : _GEN_362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_364 = 7'h22 == r_count_3_io_out ? io_r_34_b : _GEN_363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_365 = 7'h23 == r_count_3_io_out ? io_r_35_b : _GEN_364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_366 = 7'h24 == r_count_3_io_out ? io_r_36_b : _GEN_365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_367 = 7'h25 == r_count_3_io_out ? io_r_37_b : _GEN_366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_368 = 7'h26 == r_count_3_io_out ? io_r_38_b : _GEN_367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_369 = 7'h27 == r_count_3_io_out ? io_r_39_b : _GEN_368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_370 = 7'h28 == r_count_3_io_out ? io_r_40_b : _GEN_369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_371 = 7'h29 == r_count_3_io_out ? io_r_41_b : _GEN_370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_372 = 7'h2a == r_count_3_io_out ? io_r_42_b : _GEN_371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_373 = 7'h2b == r_count_3_io_out ? io_r_43_b : _GEN_372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_374 = 7'h2c == r_count_3_io_out ? io_r_44_b : _GEN_373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_375 = 7'h2d == r_count_3_io_out ? io_r_45_b : _GEN_374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_376 = 7'h2e == r_count_3_io_out ? io_r_46_b : _GEN_375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_377 = 7'h2f == r_count_3_io_out ? io_r_47_b : _GEN_376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_378 = 7'h30 == r_count_3_io_out ? io_r_48_b : _GEN_377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_379 = 7'h31 == r_count_3_io_out ? io_r_49_b : _GEN_378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_380 = 7'h32 == r_count_3_io_out ? io_r_50_b : _GEN_379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_381 = 7'h33 == r_count_3_io_out ? io_r_51_b : _GEN_380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_382 = 7'h34 == r_count_3_io_out ? io_r_52_b : _GEN_381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_383 = 7'h35 == r_count_3_io_out ? io_r_53_b : _GEN_382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_384 = 7'h36 == r_count_3_io_out ? io_r_54_b : _GEN_383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_385 = 7'h37 == r_count_3_io_out ? io_r_55_b : _GEN_384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_386 = 7'h38 == r_count_3_io_out ? io_r_56_b : _GEN_385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_387 = 7'h39 == r_count_3_io_out ? io_r_57_b : _GEN_386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_388 = 7'h3a == r_count_3_io_out ? io_r_58_b : _GEN_387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_389 = 7'h3b == r_count_3_io_out ? io_r_59_b : _GEN_388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_390 = 7'h3c == r_count_3_io_out ? io_r_60_b : _GEN_389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_391 = 7'h3d == r_count_3_io_out ? io_r_61_b : _GEN_390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_392 = 7'h3e == r_count_3_io_out ? io_r_62_b : _GEN_391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_393 = 7'h3f == r_count_3_io_out ? io_r_63_b : _GEN_392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_394 = 7'h40 == r_count_3_io_out ? io_r_64_b : _GEN_393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_395 = 7'h41 == r_count_3_io_out ? io_r_65_b : _GEN_394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_396 = 7'h42 == r_count_3_io_out ? io_r_66_b : _GEN_395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_397 = 7'h43 == r_count_3_io_out ? io_r_67_b : _GEN_396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_398 = 7'h44 == r_count_3_io_out ? io_r_68_b : _GEN_397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_399 = 7'h45 == r_count_3_io_out ? io_r_69_b : _GEN_398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_400 = 7'h46 == r_count_3_io_out ? io_r_70_b : _GEN_399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_401 = 7'h47 == r_count_3_io_out ? io_r_71_b : _GEN_400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_402 = 7'h48 == r_count_3_io_out ? io_r_72_b : _GEN_401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_403 = 7'h49 == r_count_3_io_out ? io_r_73_b : _GEN_402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_404 = 7'h4a == r_count_3_io_out ? io_r_74_b : _GEN_403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_405 = 7'h4b == r_count_3_io_out ? io_r_75_b : _GEN_404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_406 = 7'h4c == r_count_3_io_out ? io_r_76_b : _GEN_405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_407 = 7'h4d == r_count_3_io_out ? io_r_77_b : _GEN_406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_408 = 7'h4e == r_count_3_io_out ? io_r_78_b : _GEN_407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_409 = 7'h4f == r_count_3_io_out ? io_r_79_b : _GEN_408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_410 = 7'h50 == r_count_3_io_out ? io_r_80_b : _GEN_409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_411 = 7'h51 == r_count_3_io_out ? io_r_81_b : _GEN_410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_412 = 7'h52 == r_count_3_io_out ? io_r_82_b : _GEN_411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_413 = 7'h53 == r_count_3_io_out ? io_r_83_b : _GEN_412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_414 = 7'h54 == r_count_3_io_out ? io_r_84_b : _GEN_413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_415 = 7'h55 == r_count_3_io_out ? io_r_85_b : _GEN_414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_416 = 7'h56 == r_count_3_io_out ? io_r_86_b : _GEN_415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_417 = 7'h57 == r_count_3_io_out ? io_r_87_b : _GEN_416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_418 = 7'h58 == r_count_3_io_out ? io_r_88_b : _GEN_417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_419 = 7'h59 == r_count_3_io_out ? io_r_89_b : _GEN_418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_420 = 7'h5a == r_count_3_io_out ? io_r_90_b : _GEN_419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_421 = 7'h5b == r_count_3_io_out ? io_r_91_b : _GEN_420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_422 = 7'h5c == r_count_3_io_out ? io_r_92_b : _GEN_421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_423 = 7'h5d == r_count_3_io_out ? io_r_93_b : _GEN_422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_424 = 7'h5e == r_count_3_io_out ? io_r_94_b : _GEN_423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_425 = 7'h5f == r_count_3_io_out ? io_r_95_b : _GEN_424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_426 = 7'h60 == r_count_3_io_out ? io_r_96_b : _GEN_425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_427 = 7'h61 == r_count_3_io_out ? io_r_97_b : _GEN_426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_428 = 7'h62 == r_count_3_io_out ? io_r_98_b : _GEN_427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_431 = 7'h1 == r_count_4_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_432 = 7'h2 == r_count_4_io_out ? io_r_2_b : _GEN_431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_433 = 7'h3 == r_count_4_io_out ? io_r_3_b : _GEN_432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_434 = 7'h4 == r_count_4_io_out ? io_r_4_b : _GEN_433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_435 = 7'h5 == r_count_4_io_out ? io_r_5_b : _GEN_434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_436 = 7'h6 == r_count_4_io_out ? io_r_6_b : _GEN_435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_437 = 7'h7 == r_count_4_io_out ? io_r_7_b : _GEN_436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_438 = 7'h8 == r_count_4_io_out ? io_r_8_b : _GEN_437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_439 = 7'h9 == r_count_4_io_out ? io_r_9_b : _GEN_438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_440 = 7'ha == r_count_4_io_out ? io_r_10_b : _GEN_439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_441 = 7'hb == r_count_4_io_out ? io_r_11_b : _GEN_440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_442 = 7'hc == r_count_4_io_out ? io_r_12_b : _GEN_441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_443 = 7'hd == r_count_4_io_out ? io_r_13_b : _GEN_442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_444 = 7'he == r_count_4_io_out ? io_r_14_b : _GEN_443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_445 = 7'hf == r_count_4_io_out ? io_r_15_b : _GEN_444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_446 = 7'h10 == r_count_4_io_out ? io_r_16_b : _GEN_445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_447 = 7'h11 == r_count_4_io_out ? io_r_17_b : _GEN_446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_448 = 7'h12 == r_count_4_io_out ? io_r_18_b : _GEN_447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_449 = 7'h13 == r_count_4_io_out ? io_r_19_b : _GEN_448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_450 = 7'h14 == r_count_4_io_out ? io_r_20_b : _GEN_449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_451 = 7'h15 == r_count_4_io_out ? io_r_21_b : _GEN_450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_452 = 7'h16 == r_count_4_io_out ? io_r_22_b : _GEN_451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_453 = 7'h17 == r_count_4_io_out ? io_r_23_b : _GEN_452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_454 = 7'h18 == r_count_4_io_out ? io_r_24_b : _GEN_453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_455 = 7'h19 == r_count_4_io_out ? io_r_25_b : _GEN_454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_456 = 7'h1a == r_count_4_io_out ? io_r_26_b : _GEN_455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_457 = 7'h1b == r_count_4_io_out ? io_r_27_b : _GEN_456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_458 = 7'h1c == r_count_4_io_out ? io_r_28_b : _GEN_457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_459 = 7'h1d == r_count_4_io_out ? io_r_29_b : _GEN_458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_460 = 7'h1e == r_count_4_io_out ? io_r_30_b : _GEN_459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_461 = 7'h1f == r_count_4_io_out ? io_r_31_b : _GEN_460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_462 = 7'h20 == r_count_4_io_out ? io_r_32_b : _GEN_461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_463 = 7'h21 == r_count_4_io_out ? io_r_33_b : _GEN_462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_464 = 7'h22 == r_count_4_io_out ? io_r_34_b : _GEN_463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_465 = 7'h23 == r_count_4_io_out ? io_r_35_b : _GEN_464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_466 = 7'h24 == r_count_4_io_out ? io_r_36_b : _GEN_465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_467 = 7'h25 == r_count_4_io_out ? io_r_37_b : _GEN_466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_468 = 7'h26 == r_count_4_io_out ? io_r_38_b : _GEN_467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_469 = 7'h27 == r_count_4_io_out ? io_r_39_b : _GEN_468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_470 = 7'h28 == r_count_4_io_out ? io_r_40_b : _GEN_469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_471 = 7'h29 == r_count_4_io_out ? io_r_41_b : _GEN_470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_472 = 7'h2a == r_count_4_io_out ? io_r_42_b : _GEN_471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_473 = 7'h2b == r_count_4_io_out ? io_r_43_b : _GEN_472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_474 = 7'h2c == r_count_4_io_out ? io_r_44_b : _GEN_473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_475 = 7'h2d == r_count_4_io_out ? io_r_45_b : _GEN_474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_476 = 7'h2e == r_count_4_io_out ? io_r_46_b : _GEN_475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_477 = 7'h2f == r_count_4_io_out ? io_r_47_b : _GEN_476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_478 = 7'h30 == r_count_4_io_out ? io_r_48_b : _GEN_477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_479 = 7'h31 == r_count_4_io_out ? io_r_49_b : _GEN_478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_480 = 7'h32 == r_count_4_io_out ? io_r_50_b : _GEN_479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_481 = 7'h33 == r_count_4_io_out ? io_r_51_b : _GEN_480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_482 = 7'h34 == r_count_4_io_out ? io_r_52_b : _GEN_481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_483 = 7'h35 == r_count_4_io_out ? io_r_53_b : _GEN_482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_484 = 7'h36 == r_count_4_io_out ? io_r_54_b : _GEN_483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_485 = 7'h37 == r_count_4_io_out ? io_r_55_b : _GEN_484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_486 = 7'h38 == r_count_4_io_out ? io_r_56_b : _GEN_485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_487 = 7'h39 == r_count_4_io_out ? io_r_57_b : _GEN_486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_488 = 7'h3a == r_count_4_io_out ? io_r_58_b : _GEN_487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_489 = 7'h3b == r_count_4_io_out ? io_r_59_b : _GEN_488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_490 = 7'h3c == r_count_4_io_out ? io_r_60_b : _GEN_489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_491 = 7'h3d == r_count_4_io_out ? io_r_61_b : _GEN_490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_492 = 7'h3e == r_count_4_io_out ? io_r_62_b : _GEN_491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_493 = 7'h3f == r_count_4_io_out ? io_r_63_b : _GEN_492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_494 = 7'h40 == r_count_4_io_out ? io_r_64_b : _GEN_493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_495 = 7'h41 == r_count_4_io_out ? io_r_65_b : _GEN_494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_496 = 7'h42 == r_count_4_io_out ? io_r_66_b : _GEN_495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_497 = 7'h43 == r_count_4_io_out ? io_r_67_b : _GEN_496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_498 = 7'h44 == r_count_4_io_out ? io_r_68_b : _GEN_497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_499 = 7'h45 == r_count_4_io_out ? io_r_69_b : _GEN_498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_500 = 7'h46 == r_count_4_io_out ? io_r_70_b : _GEN_499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_501 = 7'h47 == r_count_4_io_out ? io_r_71_b : _GEN_500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_502 = 7'h48 == r_count_4_io_out ? io_r_72_b : _GEN_501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_503 = 7'h49 == r_count_4_io_out ? io_r_73_b : _GEN_502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_504 = 7'h4a == r_count_4_io_out ? io_r_74_b : _GEN_503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_505 = 7'h4b == r_count_4_io_out ? io_r_75_b : _GEN_504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_506 = 7'h4c == r_count_4_io_out ? io_r_76_b : _GEN_505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_507 = 7'h4d == r_count_4_io_out ? io_r_77_b : _GEN_506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_508 = 7'h4e == r_count_4_io_out ? io_r_78_b : _GEN_507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_509 = 7'h4f == r_count_4_io_out ? io_r_79_b : _GEN_508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_510 = 7'h50 == r_count_4_io_out ? io_r_80_b : _GEN_509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_511 = 7'h51 == r_count_4_io_out ? io_r_81_b : _GEN_510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_512 = 7'h52 == r_count_4_io_out ? io_r_82_b : _GEN_511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_513 = 7'h53 == r_count_4_io_out ? io_r_83_b : _GEN_512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_514 = 7'h54 == r_count_4_io_out ? io_r_84_b : _GEN_513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_515 = 7'h55 == r_count_4_io_out ? io_r_85_b : _GEN_514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_516 = 7'h56 == r_count_4_io_out ? io_r_86_b : _GEN_515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_517 = 7'h57 == r_count_4_io_out ? io_r_87_b : _GEN_516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_518 = 7'h58 == r_count_4_io_out ? io_r_88_b : _GEN_517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_519 = 7'h59 == r_count_4_io_out ? io_r_89_b : _GEN_518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_520 = 7'h5a == r_count_4_io_out ? io_r_90_b : _GEN_519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_521 = 7'h5b == r_count_4_io_out ? io_r_91_b : _GEN_520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_522 = 7'h5c == r_count_4_io_out ? io_r_92_b : _GEN_521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_523 = 7'h5d == r_count_4_io_out ? io_r_93_b : _GEN_522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_524 = 7'h5e == r_count_4_io_out ? io_r_94_b : _GEN_523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_525 = 7'h5f == r_count_4_io_out ? io_r_95_b : _GEN_524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_526 = 7'h60 == r_count_4_io_out ? io_r_96_b : _GEN_525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_527 = 7'h61 == r_count_4_io_out ? io_r_97_b : _GEN_526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_528 = 7'h62 == r_count_4_io_out ? io_r_98_b : _GEN_527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_531 = 7'h1 == r_count_5_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_532 = 7'h2 == r_count_5_io_out ? io_r_2_b : _GEN_531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_533 = 7'h3 == r_count_5_io_out ? io_r_3_b : _GEN_532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_534 = 7'h4 == r_count_5_io_out ? io_r_4_b : _GEN_533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_535 = 7'h5 == r_count_5_io_out ? io_r_5_b : _GEN_534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_536 = 7'h6 == r_count_5_io_out ? io_r_6_b : _GEN_535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_537 = 7'h7 == r_count_5_io_out ? io_r_7_b : _GEN_536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_538 = 7'h8 == r_count_5_io_out ? io_r_8_b : _GEN_537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_539 = 7'h9 == r_count_5_io_out ? io_r_9_b : _GEN_538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_540 = 7'ha == r_count_5_io_out ? io_r_10_b : _GEN_539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_541 = 7'hb == r_count_5_io_out ? io_r_11_b : _GEN_540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_542 = 7'hc == r_count_5_io_out ? io_r_12_b : _GEN_541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_543 = 7'hd == r_count_5_io_out ? io_r_13_b : _GEN_542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_544 = 7'he == r_count_5_io_out ? io_r_14_b : _GEN_543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_545 = 7'hf == r_count_5_io_out ? io_r_15_b : _GEN_544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_546 = 7'h10 == r_count_5_io_out ? io_r_16_b : _GEN_545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_547 = 7'h11 == r_count_5_io_out ? io_r_17_b : _GEN_546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_548 = 7'h12 == r_count_5_io_out ? io_r_18_b : _GEN_547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_549 = 7'h13 == r_count_5_io_out ? io_r_19_b : _GEN_548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_550 = 7'h14 == r_count_5_io_out ? io_r_20_b : _GEN_549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_551 = 7'h15 == r_count_5_io_out ? io_r_21_b : _GEN_550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_552 = 7'h16 == r_count_5_io_out ? io_r_22_b : _GEN_551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_553 = 7'h17 == r_count_5_io_out ? io_r_23_b : _GEN_552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_554 = 7'h18 == r_count_5_io_out ? io_r_24_b : _GEN_553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_555 = 7'h19 == r_count_5_io_out ? io_r_25_b : _GEN_554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_556 = 7'h1a == r_count_5_io_out ? io_r_26_b : _GEN_555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_557 = 7'h1b == r_count_5_io_out ? io_r_27_b : _GEN_556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_558 = 7'h1c == r_count_5_io_out ? io_r_28_b : _GEN_557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_559 = 7'h1d == r_count_5_io_out ? io_r_29_b : _GEN_558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_560 = 7'h1e == r_count_5_io_out ? io_r_30_b : _GEN_559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_561 = 7'h1f == r_count_5_io_out ? io_r_31_b : _GEN_560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_562 = 7'h20 == r_count_5_io_out ? io_r_32_b : _GEN_561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_563 = 7'h21 == r_count_5_io_out ? io_r_33_b : _GEN_562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_564 = 7'h22 == r_count_5_io_out ? io_r_34_b : _GEN_563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_565 = 7'h23 == r_count_5_io_out ? io_r_35_b : _GEN_564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_566 = 7'h24 == r_count_5_io_out ? io_r_36_b : _GEN_565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_567 = 7'h25 == r_count_5_io_out ? io_r_37_b : _GEN_566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_568 = 7'h26 == r_count_5_io_out ? io_r_38_b : _GEN_567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_569 = 7'h27 == r_count_5_io_out ? io_r_39_b : _GEN_568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_570 = 7'h28 == r_count_5_io_out ? io_r_40_b : _GEN_569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_571 = 7'h29 == r_count_5_io_out ? io_r_41_b : _GEN_570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_572 = 7'h2a == r_count_5_io_out ? io_r_42_b : _GEN_571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_573 = 7'h2b == r_count_5_io_out ? io_r_43_b : _GEN_572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_574 = 7'h2c == r_count_5_io_out ? io_r_44_b : _GEN_573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_575 = 7'h2d == r_count_5_io_out ? io_r_45_b : _GEN_574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_576 = 7'h2e == r_count_5_io_out ? io_r_46_b : _GEN_575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_577 = 7'h2f == r_count_5_io_out ? io_r_47_b : _GEN_576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_578 = 7'h30 == r_count_5_io_out ? io_r_48_b : _GEN_577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_579 = 7'h31 == r_count_5_io_out ? io_r_49_b : _GEN_578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_580 = 7'h32 == r_count_5_io_out ? io_r_50_b : _GEN_579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_581 = 7'h33 == r_count_5_io_out ? io_r_51_b : _GEN_580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_582 = 7'h34 == r_count_5_io_out ? io_r_52_b : _GEN_581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_583 = 7'h35 == r_count_5_io_out ? io_r_53_b : _GEN_582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_584 = 7'h36 == r_count_5_io_out ? io_r_54_b : _GEN_583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_585 = 7'h37 == r_count_5_io_out ? io_r_55_b : _GEN_584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_586 = 7'h38 == r_count_5_io_out ? io_r_56_b : _GEN_585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_587 = 7'h39 == r_count_5_io_out ? io_r_57_b : _GEN_586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_588 = 7'h3a == r_count_5_io_out ? io_r_58_b : _GEN_587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_589 = 7'h3b == r_count_5_io_out ? io_r_59_b : _GEN_588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_590 = 7'h3c == r_count_5_io_out ? io_r_60_b : _GEN_589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_591 = 7'h3d == r_count_5_io_out ? io_r_61_b : _GEN_590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_592 = 7'h3e == r_count_5_io_out ? io_r_62_b : _GEN_591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_593 = 7'h3f == r_count_5_io_out ? io_r_63_b : _GEN_592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_594 = 7'h40 == r_count_5_io_out ? io_r_64_b : _GEN_593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_595 = 7'h41 == r_count_5_io_out ? io_r_65_b : _GEN_594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_596 = 7'h42 == r_count_5_io_out ? io_r_66_b : _GEN_595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_597 = 7'h43 == r_count_5_io_out ? io_r_67_b : _GEN_596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_598 = 7'h44 == r_count_5_io_out ? io_r_68_b : _GEN_597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_599 = 7'h45 == r_count_5_io_out ? io_r_69_b : _GEN_598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_600 = 7'h46 == r_count_5_io_out ? io_r_70_b : _GEN_599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_601 = 7'h47 == r_count_5_io_out ? io_r_71_b : _GEN_600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_602 = 7'h48 == r_count_5_io_out ? io_r_72_b : _GEN_601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_603 = 7'h49 == r_count_5_io_out ? io_r_73_b : _GEN_602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_604 = 7'h4a == r_count_5_io_out ? io_r_74_b : _GEN_603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_605 = 7'h4b == r_count_5_io_out ? io_r_75_b : _GEN_604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_606 = 7'h4c == r_count_5_io_out ? io_r_76_b : _GEN_605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_607 = 7'h4d == r_count_5_io_out ? io_r_77_b : _GEN_606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_608 = 7'h4e == r_count_5_io_out ? io_r_78_b : _GEN_607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_609 = 7'h4f == r_count_5_io_out ? io_r_79_b : _GEN_608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_610 = 7'h50 == r_count_5_io_out ? io_r_80_b : _GEN_609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_611 = 7'h51 == r_count_5_io_out ? io_r_81_b : _GEN_610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_612 = 7'h52 == r_count_5_io_out ? io_r_82_b : _GEN_611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_613 = 7'h53 == r_count_5_io_out ? io_r_83_b : _GEN_612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_614 = 7'h54 == r_count_5_io_out ? io_r_84_b : _GEN_613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_615 = 7'h55 == r_count_5_io_out ? io_r_85_b : _GEN_614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_616 = 7'h56 == r_count_5_io_out ? io_r_86_b : _GEN_615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_617 = 7'h57 == r_count_5_io_out ? io_r_87_b : _GEN_616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_618 = 7'h58 == r_count_5_io_out ? io_r_88_b : _GEN_617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_619 = 7'h59 == r_count_5_io_out ? io_r_89_b : _GEN_618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_620 = 7'h5a == r_count_5_io_out ? io_r_90_b : _GEN_619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_621 = 7'h5b == r_count_5_io_out ? io_r_91_b : _GEN_620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_622 = 7'h5c == r_count_5_io_out ? io_r_92_b : _GEN_621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_623 = 7'h5d == r_count_5_io_out ? io_r_93_b : _GEN_622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_624 = 7'h5e == r_count_5_io_out ? io_r_94_b : _GEN_623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_625 = 7'h5f == r_count_5_io_out ? io_r_95_b : _GEN_624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_626 = 7'h60 == r_count_5_io_out ? io_r_96_b : _GEN_625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_627 = 7'h61 == r_count_5_io_out ? io_r_97_b : _GEN_626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_628 = 7'h62 == r_count_5_io_out ? io_r_98_b : _GEN_627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_631 = 7'h1 == r_count_6_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_632 = 7'h2 == r_count_6_io_out ? io_r_2_b : _GEN_631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_633 = 7'h3 == r_count_6_io_out ? io_r_3_b : _GEN_632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_634 = 7'h4 == r_count_6_io_out ? io_r_4_b : _GEN_633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_635 = 7'h5 == r_count_6_io_out ? io_r_5_b : _GEN_634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_636 = 7'h6 == r_count_6_io_out ? io_r_6_b : _GEN_635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_637 = 7'h7 == r_count_6_io_out ? io_r_7_b : _GEN_636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_638 = 7'h8 == r_count_6_io_out ? io_r_8_b : _GEN_637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_639 = 7'h9 == r_count_6_io_out ? io_r_9_b : _GEN_638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_640 = 7'ha == r_count_6_io_out ? io_r_10_b : _GEN_639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_641 = 7'hb == r_count_6_io_out ? io_r_11_b : _GEN_640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_642 = 7'hc == r_count_6_io_out ? io_r_12_b : _GEN_641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_643 = 7'hd == r_count_6_io_out ? io_r_13_b : _GEN_642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_644 = 7'he == r_count_6_io_out ? io_r_14_b : _GEN_643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_645 = 7'hf == r_count_6_io_out ? io_r_15_b : _GEN_644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_646 = 7'h10 == r_count_6_io_out ? io_r_16_b : _GEN_645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_647 = 7'h11 == r_count_6_io_out ? io_r_17_b : _GEN_646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_648 = 7'h12 == r_count_6_io_out ? io_r_18_b : _GEN_647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_649 = 7'h13 == r_count_6_io_out ? io_r_19_b : _GEN_648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_650 = 7'h14 == r_count_6_io_out ? io_r_20_b : _GEN_649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_651 = 7'h15 == r_count_6_io_out ? io_r_21_b : _GEN_650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_652 = 7'h16 == r_count_6_io_out ? io_r_22_b : _GEN_651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_653 = 7'h17 == r_count_6_io_out ? io_r_23_b : _GEN_652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_654 = 7'h18 == r_count_6_io_out ? io_r_24_b : _GEN_653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_655 = 7'h19 == r_count_6_io_out ? io_r_25_b : _GEN_654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_656 = 7'h1a == r_count_6_io_out ? io_r_26_b : _GEN_655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_657 = 7'h1b == r_count_6_io_out ? io_r_27_b : _GEN_656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_658 = 7'h1c == r_count_6_io_out ? io_r_28_b : _GEN_657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_659 = 7'h1d == r_count_6_io_out ? io_r_29_b : _GEN_658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_660 = 7'h1e == r_count_6_io_out ? io_r_30_b : _GEN_659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_661 = 7'h1f == r_count_6_io_out ? io_r_31_b : _GEN_660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_662 = 7'h20 == r_count_6_io_out ? io_r_32_b : _GEN_661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_663 = 7'h21 == r_count_6_io_out ? io_r_33_b : _GEN_662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_664 = 7'h22 == r_count_6_io_out ? io_r_34_b : _GEN_663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_665 = 7'h23 == r_count_6_io_out ? io_r_35_b : _GEN_664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_666 = 7'h24 == r_count_6_io_out ? io_r_36_b : _GEN_665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_667 = 7'h25 == r_count_6_io_out ? io_r_37_b : _GEN_666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_668 = 7'h26 == r_count_6_io_out ? io_r_38_b : _GEN_667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_669 = 7'h27 == r_count_6_io_out ? io_r_39_b : _GEN_668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_670 = 7'h28 == r_count_6_io_out ? io_r_40_b : _GEN_669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_671 = 7'h29 == r_count_6_io_out ? io_r_41_b : _GEN_670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_672 = 7'h2a == r_count_6_io_out ? io_r_42_b : _GEN_671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_673 = 7'h2b == r_count_6_io_out ? io_r_43_b : _GEN_672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_674 = 7'h2c == r_count_6_io_out ? io_r_44_b : _GEN_673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_675 = 7'h2d == r_count_6_io_out ? io_r_45_b : _GEN_674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_676 = 7'h2e == r_count_6_io_out ? io_r_46_b : _GEN_675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_677 = 7'h2f == r_count_6_io_out ? io_r_47_b : _GEN_676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_678 = 7'h30 == r_count_6_io_out ? io_r_48_b : _GEN_677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_679 = 7'h31 == r_count_6_io_out ? io_r_49_b : _GEN_678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_680 = 7'h32 == r_count_6_io_out ? io_r_50_b : _GEN_679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_681 = 7'h33 == r_count_6_io_out ? io_r_51_b : _GEN_680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_682 = 7'h34 == r_count_6_io_out ? io_r_52_b : _GEN_681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_683 = 7'h35 == r_count_6_io_out ? io_r_53_b : _GEN_682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_684 = 7'h36 == r_count_6_io_out ? io_r_54_b : _GEN_683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_685 = 7'h37 == r_count_6_io_out ? io_r_55_b : _GEN_684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_686 = 7'h38 == r_count_6_io_out ? io_r_56_b : _GEN_685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_687 = 7'h39 == r_count_6_io_out ? io_r_57_b : _GEN_686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_688 = 7'h3a == r_count_6_io_out ? io_r_58_b : _GEN_687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_689 = 7'h3b == r_count_6_io_out ? io_r_59_b : _GEN_688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_690 = 7'h3c == r_count_6_io_out ? io_r_60_b : _GEN_689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_691 = 7'h3d == r_count_6_io_out ? io_r_61_b : _GEN_690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_692 = 7'h3e == r_count_6_io_out ? io_r_62_b : _GEN_691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_693 = 7'h3f == r_count_6_io_out ? io_r_63_b : _GEN_692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_694 = 7'h40 == r_count_6_io_out ? io_r_64_b : _GEN_693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_695 = 7'h41 == r_count_6_io_out ? io_r_65_b : _GEN_694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_696 = 7'h42 == r_count_6_io_out ? io_r_66_b : _GEN_695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_697 = 7'h43 == r_count_6_io_out ? io_r_67_b : _GEN_696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_698 = 7'h44 == r_count_6_io_out ? io_r_68_b : _GEN_697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_699 = 7'h45 == r_count_6_io_out ? io_r_69_b : _GEN_698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_700 = 7'h46 == r_count_6_io_out ? io_r_70_b : _GEN_699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_701 = 7'h47 == r_count_6_io_out ? io_r_71_b : _GEN_700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_702 = 7'h48 == r_count_6_io_out ? io_r_72_b : _GEN_701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_703 = 7'h49 == r_count_6_io_out ? io_r_73_b : _GEN_702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_704 = 7'h4a == r_count_6_io_out ? io_r_74_b : _GEN_703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_705 = 7'h4b == r_count_6_io_out ? io_r_75_b : _GEN_704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_706 = 7'h4c == r_count_6_io_out ? io_r_76_b : _GEN_705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_707 = 7'h4d == r_count_6_io_out ? io_r_77_b : _GEN_706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_708 = 7'h4e == r_count_6_io_out ? io_r_78_b : _GEN_707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_709 = 7'h4f == r_count_6_io_out ? io_r_79_b : _GEN_708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_710 = 7'h50 == r_count_6_io_out ? io_r_80_b : _GEN_709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_711 = 7'h51 == r_count_6_io_out ? io_r_81_b : _GEN_710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_712 = 7'h52 == r_count_6_io_out ? io_r_82_b : _GEN_711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_713 = 7'h53 == r_count_6_io_out ? io_r_83_b : _GEN_712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_714 = 7'h54 == r_count_6_io_out ? io_r_84_b : _GEN_713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_715 = 7'h55 == r_count_6_io_out ? io_r_85_b : _GEN_714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_716 = 7'h56 == r_count_6_io_out ? io_r_86_b : _GEN_715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_717 = 7'h57 == r_count_6_io_out ? io_r_87_b : _GEN_716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_718 = 7'h58 == r_count_6_io_out ? io_r_88_b : _GEN_717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_719 = 7'h59 == r_count_6_io_out ? io_r_89_b : _GEN_718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_720 = 7'h5a == r_count_6_io_out ? io_r_90_b : _GEN_719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_721 = 7'h5b == r_count_6_io_out ? io_r_91_b : _GEN_720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_722 = 7'h5c == r_count_6_io_out ? io_r_92_b : _GEN_721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_723 = 7'h5d == r_count_6_io_out ? io_r_93_b : _GEN_722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_724 = 7'h5e == r_count_6_io_out ? io_r_94_b : _GEN_723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_725 = 7'h5f == r_count_6_io_out ? io_r_95_b : _GEN_724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_726 = 7'h60 == r_count_6_io_out ? io_r_96_b : _GEN_725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_727 = 7'h61 == r_count_6_io_out ? io_r_97_b : _GEN_726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_728 = 7'h62 == r_count_6_io_out ? io_r_98_b : _GEN_727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_731 = 7'h1 == r_count_7_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_732 = 7'h2 == r_count_7_io_out ? io_r_2_b : _GEN_731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_733 = 7'h3 == r_count_7_io_out ? io_r_3_b : _GEN_732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_734 = 7'h4 == r_count_7_io_out ? io_r_4_b : _GEN_733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_735 = 7'h5 == r_count_7_io_out ? io_r_5_b : _GEN_734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_736 = 7'h6 == r_count_7_io_out ? io_r_6_b : _GEN_735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_737 = 7'h7 == r_count_7_io_out ? io_r_7_b : _GEN_736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_738 = 7'h8 == r_count_7_io_out ? io_r_8_b : _GEN_737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_739 = 7'h9 == r_count_7_io_out ? io_r_9_b : _GEN_738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_740 = 7'ha == r_count_7_io_out ? io_r_10_b : _GEN_739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_741 = 7'hb == r_count_7_io_out ? io_r_11_b : _GEN_740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_742 = 7'hc == r_count_7_io_out ? io_r_12_b : _GEN_741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_743 = 7'hd == r_count_7_io_out ? io_r_13_b : _GEN_742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_744 = 7'he == r_count_7_io_out ? io_r_14_b : _GEN_743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_745 = 7'hf == r_count_7_io_out ? io_r_15_b : _GEN_744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_746 = 7'h10 == r_count_7_io_out ? io_r_16_b : _GEN_745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_747 = 7'h11 == r_count_7_io_out ? io_r_17_b : _GEN_746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_748 = 7'h12 == r_count_7_io_out ? io_r_18_b : _GEN_747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_749 = 7'h13 == r_count_7_io_out ? io_r_19_b : _GEN_748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_750 = 7'h14 == r_count_7_io_out ? io_r_20_b : _GEN_749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_751 = 7'h15 == r_count_7_io_out ? io_r_21_b : _GEN_750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_752 = 7'h16 == r_count_7_io_out ? io_r_22_b : _GEN_751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_753 = 7'h17 == r_count_7_io_out ? io_r_23_b : _GEN_752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_754 = 7'h18 == r_count_7_io_out ? io_r_24_b : _GEN_753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_755 = 7'h19 == r_count_7_io_out ? io_r_25_b : _GEN_754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_756 = 7'h1a == r_count_7_io_out ? io_r_26_b : _GEN_755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_757 = 7'h1b == r_count_7_io_out ? io_r_27_b : _GEN_756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_758 = 7'h1c == r_count_7_io_out ? io_r_28_b : _GEN_757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_759 = 7'h1d == r_count_7_io_out ? io_r_29_b : _GEN_758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_760 = 7'h1e == r_count_7_io_out ? io_r_30_b : _GEN_759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_761 = 7'h1f == r_count_7_io_out ? io_r_31_b : _GEN_760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_762 = 7'h20 == r_count_7_io_out ? io_r_32_b : _GEN_761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_763 = 7'h21 == r_count_7_io_out ? io_r_33_b : _GEN_762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_764 = 7'h22 == r_count_7_io_out ? io_r_34_b : _GEN_763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_765 = 7'h23 == r_count_7_io_out ? io_r_35_b : _GEN_764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_766 = 7'h24 == r_count_7_io_out ? io_r_36_b : _GEN_765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_767 = 7'h25 == r_count_7_io_out ? io_r_37_b : _GEN_766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_768 = 7'h26 == r_count_7_io_out ? io_r_38_b : _GEN_767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_769 = 7'h27 == r_count_7_io_out ? io_r_39_b : _GEN_768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_770 = 7'h28 == r_count_7_io_out ? io_r_40_b : _GEN_769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_771 = 7'h29 == r_count_7_io_out ? io_r_41_b : _GEN_770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_772 = 7'h2a == r_count_7_io_out ? io_r_42_b : _GEN_771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_773 = 7'h2b == r_count_7_io_out ? io_r_43_b : _GEN_772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_774 = 7'h2c == r_count_7_io_out ? io_r_44_b : _GEN_773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_775 = 7'h2d == r_count_7_io_out ? io_r_45_b : _GEN_774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_776 = 7'h2e == r_count_7_io_out ? io_r_46_b : _GEN_775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_777 = 7'h2f == r_count_7_io_out ? io_r_47_b : _GEN_776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_778 = 7'h30 == r_count_7_io_out ? io_r_48_b : _GEN_777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_779 = 7'h31 == r_count_7_io_out ? io_r_49_b : _GEN_778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_780 = 7'h32 == r_count_7_io_out ? io_r_50_b : _GEN_779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_781 = 7'h33 == r_count_7_io_out ? io_r_51_b : _GEN_780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_782 = 7'h34 == r_count_7_io_out ? io_r_52_b : _GEN_781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_783 = 7'h35 == r_count_7_io_out ? io_r_53_b : _GEN_782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_784 = 7'h36 == r_count_7_io_out ? io_r_54_b : _GEN_783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_785 = 7'h37 == r_count_7_io_out ? io_r_55_b : _GEN_784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_786 = 7'h38 == r_count_7_io_out ? io_r_56_b : _GEN_785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_787 = 7'h39 == r_count_7_io_out ? io_r_57_b : _GEN_786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_788 = 7'h3a == r_count_7_io_out ? io_r_58_b : _GEN_787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_789 = 7'h3b == r_count_7_io_out ? io_r_59_b : _GEN_788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_790 = 7'h3c == r_count_7_io_out ? io_r_60_b : _GEN_789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_791 = 7'h3d == r_count_7_io_out ? io_r_61_b : _GEN_790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_792 = 7'h3e == r_count_7_io_out ? io_r_62_b : _GEN_791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_793 = 7'h3f == r_count_7_io_out ? io_r_63_b : _GEN_792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_794 = 7'h40 == r_count_7_io_out ? io_r_64_b : _GEN_793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_795 = 7'h41 == r_count_7_io_out ? io_r_65_b : _GEN_794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_796 = 7'h42 == r_count_7_io_out ? io_r_66_b : _GEN_795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_797 = 7'h43 == r_count_7_io_out ? io_r_67_b : _GEN_796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_798 = 7'h44 == r_count_7_io_out ? io_r_68_b : _GEN_797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_799 = 7'h45 == r_count_7_io_out ? io_r_69_b : _GEN_798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_800 = 7'h46 == r_count_7_io_out ? io_r_70_b : _GEN_799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_801 = 7'h47 == r_count_7_io_out ? io_r_71_b : _GEN_800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_802 = 7'h48 == r_count_7_io_out ? io_r_72_b : _GEN_801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_803 = 7'h49 == r_count_7_io_out ? io_r_73_b : _GEN_802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_804 = 7'h4a == r_count_7_io_out ? io_r_74_b : _GEN_803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_805 = 7'h4b == r_count_7_io_out ? io_r_75_b : _GEN_804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_806 = 7'h4c == r_count_7_io_out ? io_r_76_b : _GEN_805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_807 = 7'h4d == r_count_7_io_out ? io_r_77_b : _GEN_806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_808 = 7'h4e == r_count_7_io_out ? io_r_78_b : _GEN_807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_809 = 7'h4f == r_count_7_io_out ? io_r_79_b : _GEN_808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_810 = 7'h50 == r_count_7_io_out ? io_r_80_b : _GEN_809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_811 = 7'h51 == r_count_7_io_out ? io_r_81_b : _GEN_810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_812 = 7'h52 == r_count_7_io_out ? io_r_82_b : _GEN_811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_813 = 7'h53 == r_count_7_io_out ? io_r_83_b : _GEN_812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_814 = 7'h54 == r_count_7_io_out ? io_r_84_b : _GEN_813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_815 = 7'h55 == r_count_7_io_out ? io_r_85_b : _GEN_814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_816 = 7'h56 == r_count_7_io_out ? io_r_86_b : _GEN_815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_817 = 7'h57 == r_count_7_io_out ? io_r_87_b : _GEN_816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_818 = 7'h58 == r_count_7_io_out ? io_r_88_b : _GEN_817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_819 = 7'h59 == r_count_7_io_out ? io_r_89_b : _GEN_818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_820 = 7'h5a == r_count_7_io_out ? io_r_90_b : _GEN_819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_821 = 7'h5b == r_count_7_io_out ? io_r_91_b : _GEN_820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_822 = 7'h5c == r_count_7_io_out ? io_r_92_b : _GEN_821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_823 = 7'h5d == r_count_7_io_out ? io_r_93_b : _GEN_822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_824 = 7'h5e == r_count_7_io_out ? io_r_94_b : _GEN_823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_825 = 7'h5f == r_count_7_io_out ? io_r_95_b : _GEN_824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_826 = 7'h60 == r_count_7_io_out ? io_r_96_b : _GEN_825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_827 = 7'h61 == r_count_7_io_out ? io_r_97_b : _GEN_826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_828 = 7'h62 == r_count_7_io_out ? io_r_98_b : _GEN_827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_831 = 7'h1 == r_count_8_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_832 = 7'h2 == r_count_8_io_out ? io_r_2_b : _GEN_831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_833 = 7'h3 == r_count_8_io_out ? io_r_3_b : _GEN_832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_834 = 7'h4 == r_count_8_io_out ? io_r_4_b : _GEN_833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_835 = 7'h5 == r_count_8_io_out ? io_r_5_b : _GEN_834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_836 = 7'h6 == r_count_8_io_out ? io_r_6_b : _GEN_835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_837 = 7'h7 == r_count_8_io_out ? io_r_7_b : _GEN_836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_838 = 7'h8 == r_count_8_io_out ? io_r_8_b : _GEN_837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_839 = 7'h9 == r_count_8_io_out ? io_r_9_b : _GEN_838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_840 = 7'ha == r_count_8_io_out ? io_r_10_b : _GEN_839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_841 = 7'hb == r_count_8_io_out ? io_r_11_b : _GEN_840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_842 = 7'hc == r_count_8_io_out ? io_r_12_b : _GEN_841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_843 = 7'hd == r_count_8_io_out ? io_r_13_b : _GEN_842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_844 = 7'he == r_count_8_io_out ? io_r_14_b : _GEN_843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_845 = 7'hf == r_count_8_io_out ? io_r_15_b : _GEN_844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_846 = 7'h10 == r_count_8_io_out ? io_r_16_b : _GEN_845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_847 = 7'h11 == r_count_8_io_out ? io_r_17_b : _GEN_846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_848 = 7'h12 == r_count_8_io_out ? io_r_18_b : _GEN_847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_849 = 7'h13 == r_count_8_io_out ? io_r_19_b : _GEN_848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_850 = 7'h14 == r_count_8_io_out ? io_r_20_b : _GEN_849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_851 = 7'h15 == r_count_8_io_out ? io_r_21_b : _GEN_850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_852 = 7'h16 == r_count_8_io_out ? io_r_22_b : _GEN_851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_853 = 7'h17 == r_count_8_io_out ? io_r_23_b : _GEN_852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_854 = 7'h18 == r_count_8_io_out ? io_r_24_b : _GEN_853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_855 = 7'h19 == r_count_8_io_out ? io_r_25_b : _GEN_854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_856 = 7'h1a == r_count_8_io_out ? io_r_26_b : _GEN_855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_857 = 7'h1b == r_count_8_io_out ? io_r_27_b : _GEN_856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_858 = 7'h1c == r_count_8_io_out ? io_r_28_b : _GEN_857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_859 = 7'h1d == r_count_8_io_out ? io_r_29_b : _GEN_858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_860 = 7'h1e == r_count_8_io_out ? io_r_30_b : _GEN_859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_861 = 7'h1f == r_count_8_io_out ? io_r_31_b : _GEN_860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_862 = 7'h20 == r_count_8_io_out ? io_r_32_b : _GEN_861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_863 = 7'h21 == r_count_8_io_out ? io_r_33_b : _GEN_862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_864 = 7'h22 == r_count_8_io_out ? io_r_34_b : _GEN_863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_865 = 7'h23 == r_count_8_io_out ? io_r_35_b : _GEN_864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_866 = 7'h24 == r_count_8_io_out ? io_r_36_b : _GEN_865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_867 = 7'h25 == r_count_8_io_out ? io_r_37_b : _GEN_866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_868 = 7'h26 == r_count_8_io_out ? io_r_38_b : _GEN_867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_869 = 7'h27 == r_count_8_io_out ? io_r_39_b : _GEN_868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_870 = 7'h28 == r_count_8_io_out ? io_r_40_b : _GEN_869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_871 = 7'h29 == r_count_8_io_out ? io_r_41_b : _GEN_870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_872 = 7'h2a == r_count_8_io_out ? io_r_42_b : _GEN_871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_873 = 7'h2b == r_count_8_io_out ? io_r_43_b : _GEN_872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_874 = 7'h2c == r_count_8_io_out ? io_r_44_b : _GEN_873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_875 = 7'h2d == r_count_8_io_out ? io_r_45_b : _GEN_874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_876 = 7'h2e == r_count_8_io_out ? io_r_46_b : _GEN_875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_877 = 7'h2f == r_count_8_io_out ? io_r_47_b : _GEN_876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_878 = 7'h30 == r_count_8_io_out ? io_r_48_b : _GEN_877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_879 = 7'h31 == r_count_8_io_out ? io_r_49_b : _GEN_878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_880 = 7'h32 == r_count_8_io_out ? io_r_50_b : _GEN_879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_881 = 7'h33 == r_count_8_io_out ? io_r_51_b : _GEN_880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_882 = 7'h34 == r_count_8_io_out ? io_r_52_b : _GEN_881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_883 = 7'h35 == r_count_8_io_out ? io_r_53_b : _GEN_882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_884 = 7'h36 == r_count_8_io_out ? io_r_54_b : _GEN_883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_885 = 7'h37 == r_count_8_io_out ? io_r_55_b : _GEN_884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_886 = 7'h38 == r_count_8_io_out ? io_r_56_b : _GEN_885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_887 = 7'h39 == r_count_8_io_out ? io_r_57_b : _GEN_886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_888 = 7'h3a == r_count_8_io_out ? io_r_58_b : _GEN_887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_889 = 7'h3b == r_count_8_io_out ? io_r_59_b : _GEN_888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_890 = 7'h3c == r_count_8_io_out ? io_r_60_b : _GEN_889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_891 = 7'h3d == r_count_8_io_out ? io_r_61_b : _GEN_890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_892 = 7'h3e == r_count_8_io_out ? io_r_62_b : _GEN_891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_893 = 7'h3f == r_count_8_io_out ? io_r_63_b : _GEN_892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_894 = 7'h40 == r_count_8_io_out ? io_r_64_b : _GEN_893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_895 = 7'h41 == r_count_8_io_out ? io_r_65_b : _GEN_894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_896 = 7'h42 == r_count_8_io_out ? io_r_66_b : _GEN_895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_897 = 7'h43 == r_count_8_io_out ? io_r_67_b : _GEN_896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_898 = 7'h44 == r_count_8_io_out ? io_r_68_b : _GEN_897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_899 = 7'h45 == r_count_8_io_out ? io_r_69_b : _GEN_898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_900 = 7'h46 == r_count_8_io_out ? io_r_70_b : _GEN_899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_901 = 7'h47 == r_count_8_io_out ? io_r_71_b : _GEN_900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_902 = 7'h48 == r_count_8_io_out ? io_r_72_b : _GEN_901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_903 = 7'h49 == r_count_8_io_out ? io_r_73_b : _GEN_902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_904 = 7'h4a == r_count_8_io_out ? io_r_74_b : _GEN_903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_905 = 7'h4b == r_count_8_io_out ? io_r_75_b : _GEN_904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_906 = 7'h4c == r_count_8_io_out ? io_r_76_b : _GEN_905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_907 = 7'h4d == r_count_8_io_out ? io_r_77_b : _GEN_906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_908 = 7'h4e == r_count_8_io_out ? io_r_78_b : _GEN_907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_909 = 7'h4f == r_count_8_io_out ? io_r_79_b : _GEN_908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_910 = 7'h50 == r_count_8_io_out ? io_r_80_b : _GEN_909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_911 = 7'h51 == r_count_8_io_out ? io_r_81_b : _GEN_910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_912 = 7'h52 == r_count_8_io_out ? io_r_82_b : _GEN_911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_913 = 7'h53 == r_count_8_io_out ? io_r_83_b : _GEN_912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_914 = 7'h54 == r_count_8_io_out ? io_r_84_b : _GEN_913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_915 = 7'h55 == r_count_8_io_out ? io_r_85_b : _GEN_914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_916 = 7'h56 == r_count_8_io_out ? io_r_86_b : _GEN_915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_917 = 7'h57 == r_count_8_io_out ? io_r_87_b : _GEN_916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_918 = 7'h58 == r_count_8_io_out ? io_r_88_b : _GEN_917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_919 = 7'h59 == r_count_8_io_out ? io_r_89_b : _GEN_918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_920 = 7'h5a == r_count_8_io_out ? io_r_90_b : _GEN_919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_921 = 7'h5b == r_count_8_io_out ? io_r_91_b : _GEN_920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_922 = 7'h5c == r_count_8_io_out ? io_r_92_b : _GEN_921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_923 = 7'h5d == r_count_8_io_out ? io_r_93_b : _GEN_922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_924 = 7'h5e == r_count_8_io_out ? io_r_94_b : _GEN_923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_925 = 7'h5f == r_count_8_io_out ? io_r_95_b : _GEN_924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_926 = 7'h60 == r_count_8_io_out ? io_r_96_b : _GEN_925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_927 = 7'h61 == r_count_8_io_out ? io_r_97_b : _GEN_926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_928 = 7'h62 == r_count_8_io_out ? io_r_98_b : _GEN_927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_931 = 7'h1 == r_count_9_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_932 = 7'h2 == r_count_9_io_out ? io_r_2_b : _GEN_931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_933 = 7'h3 == r_count_9_io_out ? io_r_3_b : _GEN_932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_934 = 7'h4 == r_count_9_io_out ? io_r_4_b : _GEN_933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_935 = 7'h5 == r_count_9_io_out ? io_r_5_b : _GEN_934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_936 = 7'h6 == r_count_9_io_out ? io_r_6_b : _GEN_935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_937 = 7'h7 == r_count_9_io_out ? io_r_7_b : _GEN_936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_938 = 7'h8 == r_count_9_io_out ? io_r_8_b : _GEN_937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_939 = 7'h9 == r_count_9_io_out ? io_r_9_b : _GEN_938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_940 = 7'ha == r_count_9_io_out ? io_r_10_b : _GEN_939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_941 = 7'hb == r_count_9_io_out ? io_r_11_b : _GEN_940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_942 = 7'hc == r_count_9_io_out ? io_r_12_b : _GEN_941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_943 = 7'hd == r_count_9_io_out ? io_r_13_b : _GEN_942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_944 = 7'he == r_count_9_io_out ? io_r_14_b : _GEN_943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_945 = 7'hf == r_count_9_io_out ? io_r_15_b : _GEN_944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_946 = 7'h10 == r_count_9_io_out ? io_r_16_b : _GEN_945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_947 = 7'h11 == r_count_9_io_out ? io_r_17_b : _GEN_946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_948 = 7'h12 == r_count_9_io_out ? io_r_18_b : _GEN_947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_949 = 7'h13 == r_count_9_io_out ? io_r_19_b : _GEN_948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_950 = 7'h14 == r_count_9_io_out ? io_r_20_b : _GEN_949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_951 = 7'h15 == r_count_9_io_out ? io_r_21_b : _GEN_950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_952 = 7'h16 == r_count_9_io_out ? io_r_22_b : _GEN_951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_953 = 7'h17 == r_count_9_io_out ? io_r_23_b : _GEN_952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_954 = 7'h18 == r_count_9_io_out ? io_r_24_b : _GEN_953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_955 = 7'h19 == r_count_9_io_out ? io_r_25_b : _GEN_954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_956 = 7'h1a == r_count_9_io_out ? io_r_26_b : _GEN_955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_957 = 7'h1b == r_count_9_io_out ? io_r_27_b : _GEN_956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_958 = 7'h1c == r_count_9_io_out ? io_r_28_b : _GEN_957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_959 = 7'h1d == r_count_9_io_out ? io_r_29_b : _GEN_958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_960 = 7'h1e == r_count_9_io_out ? io_r_30_b : _GEN_959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_961 = 7'h1f == r_count_9_io_out ? io_r_31_b : _GEN_960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_962 = 7'h20 == r_count_9_io_out ? io_r_32_b : _GEN_961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_963 = 7'h21 == r_count_9_io_out ? io_r_33_b : _GEN_962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_964 = 7'h22 == r_count_9_io_out ? io_r_34_b : _GEN_963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_965 = 7'h23 == r_count_9_io_out ? io_r_35_b : _GEN_964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_966 = 7'h24 == r_count_9_io_out ? io_r_36_b : _GEN_965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_967 = 7'h25 == r_count_9_io_out ? io_r_37_b : _GEN_966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_968 = 7'h26 == r_count_9_io_out ? io_r_38_b : _GEN_967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_969 = 7'h27 == r_count_9_io_out ? io_r_39_b : _GEN_968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_970 = 7'h28 == r_count_9_io_out ? io_r_40_b : _GEN_969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_971 = 7'h29 == r_count_9_io_out ? io_r_41_b : _GEN_970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_972 = 7'h2a == r_count_9_io_out ? io_r_42_b : _GEN_971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_973 = 7'h2b == r_count_9_io_out ? io_r_43_b : _GEN_972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_974 = 7'h2c == r_count_9_io_out ? io_r_44_b : _GEN_973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_975 = 7'h2d == r_count_9_io_out ? io_r_45_b : _GEN_974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_976 = 7'h2e == r_count_9_io_out ? io_r_46_b : _GEN_975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_977 = 7'h2f == r_count_9_io_out ? io_r_47_b : _GEN_976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_978 = 7'h30 == r_count_9_io_out ? io_r_48_b : _GEN_977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_979 = 7'h31 == r_count_9_io_out ? io_r_49_b : _GEN_978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_980 = 7'h32 == r_count_9_io_out ? io_r_50_b : _GEN_979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_981 = 7'h33 == r_count_9_io_out ? io_r_51_b : _GEN_980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_982 = 7'h34 == r_count_9_io_out ? io_r_52_b : _GEN_981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_983 = 7'h35 == r_count_9_io_out ? io_r_53_b : _GEN_982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_984 = 7'h36 == r_count_9_io_out ? io_r_54_b : _GEN_983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_985 = 7'h37 == r_count_9_io_out ? io_r_55_b : _GEN_984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_986 = 7'h38 == r_count_9_io_out ? io_r_56_b : _GEN_985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_987 = 7'h39 == r_count_9_io_out ? io_r_57_b : _GEN_986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_988 = 7'h3a == r_count_9_io_out ? io_r_58_b : _GEN_987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_989 = 7'h3b == r_count_9_io_out ? io_r_59_b : _GEN_988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_990 = 7'h3c == r_count_9_io_out ? io_r_60_b : _GEN_989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_991 = 7'h3d == r_count_9_io_out ? io_r_61_b : _GEN_990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_992 = 7'h3e == r_count_9_io_out ? io_r_62_b : _GEN_991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_993 = 7'h3f == r_count_9_io_out ? io_r_63_b : _GEN_992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_994 = 7'h40 == r_count_9_io_out ? io_r_64_b : _GEN_993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_995 = 7'h41 == r_count_9_io_out ? io_r_65_b : _GEN_994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_996 = 7'h42 == r_count_9_io_out ? io_r_66_b : _GEN_995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_997 = 7'h43 == r_count_9_io_out ? io_r_67_b : _GEN_996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_998 = 7'h44 == r_count_9_io_out ? io_r_68_b : _GEN_997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_999 = 7'h45 == r_count_9_io_out ? io_r_69_b : _GEN_998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1000 = 7'h46 == r_count_9_io_out ? io_r_70_b : _GEN_999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1001 = 7'h47 == r_count_9_io_out ? io_r_71_b : _GEN_1000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1002 = 7'h48 == r_count_9_io_out ? io_r_72_b : _GEN_1001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1003 = 7'h49 == r_count_9_io_out ? io_r_73_b : _GEN_1002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1004 = 7'h4a == r_count_9_io_out ? io_r_74_b : _GEN_1003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1005 = 7'h4b == r_count_9_io_out ? io_r_75_b : _GEN_1004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1006 = 7'h4c == r_count_9_io_out ? io_r_76_b : _GEN_1005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1007 = 7'h4d == r_count_9_io_out ? io_r_77_b : _GEN_1006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1008 = 7'h4e == r_count_9_io_out ? io_r_78_b : _GEN_1007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1009 = 7'h4f == r_count_9_io_out ? io_r_79_b : _GEN_1008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1010 = 7'h50 == r_count_9_io_out ? io_r_80_b : _GEN_1009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1011 = 7'h51 == r_count_9_io_out ? io_r_81_b : _GEN_1010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1012 = 7'h52 == r_count_9_io_out ? io_r_82_b : _GEN_1011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1013 = 7'h53 == r_count_9_io_out ? io_r_83_b : _GEN_1012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1014 = 7'h54 == r_count_9_io_out ? io_r_84_b : _GEN_1013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1015 = 7'h55 == r_count_9_io_out ? io_r_85_b : _GEN_1014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1016 = 7'h56 == r_count_9_io_out ? io_r_86_b : _GEN_1015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1017 = 7'h57 == r_count_9_io_out ? io_r_87_b : _GEN_1016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1018 = 7'h58 == r_count_9_io_out ? io_r_88_b : _GEN_1017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1019 = 7'h59 == r_count_9_io_out ? io_r_89_b : _GEN_1018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1020 = 7'h5a == r_count_9_io_out ? io_r_90_b : _GEN_1019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1021 = 7'h5b == r_count_9_io_out ? io_r_91_b : _GEN_1020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1022 = 7'h5c == r_count_9_io_out ? io_r_92_b : _GEN_1021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1023 = 7'h5d == r_count_9_io_out ? io_r_93_b : _GEN_1022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1024 = 7'h5e == r_count_9_io_out ? io_r_94_b : _GEN_1023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1025 = 7'h5f == r_count_9_io_out ? io_r_95_b : _GEN_1024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1026 = 7'h60 == r_count_9_io_out ? io_r_96_b : _GEN_1025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1027 = 7'h61 == r_count_9_io_out ? io_r_97_b : _GEN_1026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1028 = 7'h62 == r_count_9_io_out ? io_r_98_b : _GEN_1027; // @[SWChisel.scala 221:{19,19}]
  SWCell array_0 ( // @[SWChisel.scala 170:39]
    .io_q(array_0_io_q),
    .io_r(array_0_io_r),
    .io_e_i(array_0_io_e_i),
    .io_f_i(array_0_io_f_i),
    .io_ve_i(array_0_io_ve_i),
    .io_vf_i(array_0_io_vf_i),
    .io_vv_i(array_0_io_vv_i),
    .io_e_o(array_0_io_e_o),
    .io_f_o(array_0_io_f_o),
    .io_v_o(array_0_io_v_o)
  );
  SWCell array_1 ( // @[SWChisel.scala 170:39]
    .io_q(array_1_io_q),
    .io_r(array_1_io_r),
    .io_e_i(array_1_io_e_i),
    .io_f_i(array_1_io_f_i),
    .io_ve_i(array_1_io_ve_i),
    .io_vf_i(array_1_io_vf_i),
    .io_vv_i(array_1_io_vv_i),
    .io_e_o(array_1_io_e_o),
    .io_f_o(array_1_io_f_o),
    .io_v_o(array_1_io_v_o)
  );
  SWCell array_2 ( // @[SWChisel.scala 170:39]
    .io_q(array_2_io_q),
    .io_r(array_2_io_r),
    .io_e_i(array_2_io_e_i),
    .io_f_i(array_2_io_f_i),
    .io_ve_i(array_2_io_ve_i),
    .io_vf_i(array_2_io_vf_i),
    .io_vv_i(array_2_io_vv_i),
    .io_e_o(array_2_io_e_o),
    .io_f_o(array_2_io_f_o),
    .io_v_o(array_2_io_v_o)
  );
  SWCell array_3 ( // @[SWChisel.scala 170:39]
    .io_q(array_3_io_q),
    .io_r(array_3_io_r),
    .io_e_i(array_3_io_e_i),
    .io_f_i(array_3_io_f_i),
    .io_ve_i(array_3_io_ve_i),
    .io_vf_i(array_3_io_vf_i),
    .io_vv_i(array_3_io_vv_i),
    .io_e_o(array_3_io_e_o),
    .io_f_o(array_3_io_f_o),
    .io_v_o(array_3_io_v_o)
  );
  SWCell array_4 ( // @[SWChisel.scala 170:39]
    .io_q(array_4_io_q),
    .io_r(array_4_io_r),
    .io_e_i(array_4_io_e_i),
    .io_f_i(array_4_io_f_i),
    .io_ve_i(array_4_io_ve_i),
    .io_vf_i(array_4_io_vf_i),
    .io_vv_i(array_4_io_vv_i),
    .io_e_o(array_4_io_e_o),
    .io_f_o(array_4_io_f_o),
    .io_v_o(array_4_io_v_o)
  );
  SWCell array_5 ( // @[SWChisel.scala 170:39]
    .io_q(array_5_io_q),
    .io_r(array_5_io_r),
    .io_e_i(array_5_io_e_i),
    .io_f_i(array_5_io_f_i),
    .io_ve_i(array_5_io_ve_i),
    .io_vf_i(array_5_io_vf_i),
    .io_vv_i(array_5_io_vv_i),
    .io_e_o(array_5_io_e_o),
    .io_f_o(array_5_io_f_o),
    .io_v_o(array_5_io_v_o)
  );
  SWCell array_6 ( // @[SWChisel.scala 170:39]
    .io_q(array_6_io_q),
    .io_r(array_6_io_r),
    .io_e_i(array_6_io_e_i),
    .io_f_i(array_6_io_f_i),
    .io_ve_i(array_6_io_ve_i),
    .io_vf_i(array_6_io_vf_i),
    .io_vv_i(array_6_io_vv_i),
    .io_e_o(array_6_io_e_o),
    .io_f_o(array_6_io_f_o),
    .io_v_o(array_6_io_v_o)
  );
  SWCell array_7 ( // @[SWChisel.scala 170:39]
    .io_q(array_7_io_q),
    .io_r(array_7_io_r),
    .io_e_i(array_7_io_e_i),
    .io_f_i(array_7_io_f_i),
    .io_ve_i(array_7_io_ve_i),
    .io_vf_i(array_7_io_vf_i),
    .io_vv_i(array_7_io_vv_i),
    .io_e_o(array_7_io_e_o),
    .io_f_o(array_7_io_f_o),
    .io_v_o(array_7_io_v_o)
  );
  SWCell array_8 ( // @[SWChisel.scala 170:39]
    .io_q(array_8_io_q),
    .io_r(array_8_io_r),
    .io_e_i(array_8_io_e_i),
    .io_f_i(array_8_io_f_i),
    .io_ve_i(array_8_io_ve_i),
    .io_vf_i(array_8_io_vf_i),
    .io_vv_i(array_8_io_vv_i),
    .io_e_o(array_8_io_e_o),
    .io_f_o(array_8_io_f_o),
    .io_v_o(array_8_io_v_o)
  );
  SWCell array_9 ( // @[SWChisel.scala 170:39]
    .io_q(array_9_io_q),
    .io_r(array_9_io_r),
    .io_e_i(array_9_io_e_i),
    .io_f_i(array_9_io_f_i),
    .io_ve_i(array_9_io_ve_i),
    .io_vf_i(array_9_io_vf_i),
    .io_vv_i(array_9_io_vv_i),
    .io_e_o(array_9_io_e_o),
    .io_f_o(array_9_io_f_o),
    .io_v_o(array_9_io_v_o)
  );
  MyCounter r_count_0 ( // @[SWChisel.scala 171:41]
    .clock(r_count_0_clock),
    .reset(r_count_0_reset),
    .io_en(r_count_0_io_en),
    .io_out(r_count_0_io_out)
  );
  MyCounter r_count_1 ( // @[SWChisel.scala 171:41]
    .clock(r_count_1_clock),
    .reset(r_count_1_reset),
    .io_en(r_count_1_io_en),
    .io_out(r_count_1_io_out)
  );
  MyCounter r_count_2 ( // @[SWChisel.scala 171:41]
    .clock(r_count_2_clock),
    .reset(r_count_2_reset),
    .io_en(r_count_2_io_en),
    .io_out(r_count_2_io_out)
  );
  MyCounter r_count_3 ( // @[SWChisel.scala 171:41]
    .clock(r_count_3_clock),
    .reset(r_count_3_reset),
    .io_en(r_count_3_io_en),
    .io_out(r_count_3_io_out)
  );
  MyCounter r_count_4 ( // @[SWChisel.scala 171:41]
    .clock(r_count_4_clock),
    .reset(r_count_4_reset),
    .io_en(r_count_4_io_en),
    .io_out(r_count_4_io_out)
  );
  MyCounter r_count_5 ( // @[SWChisel.scala 171:41]
    .clock(r_count_5_clock),
    .reset(r_count_5_reset),
    .io_en(r_count_5_io_en),
    .io_out(r_count_5_io_out)
  );
  MyCounter r_count_6 ( // @[SWChisel.scala 171:41]
    .clock(r_count_6_clock),
    .reset(r_count_6_reset),
    .io_en(r_count_6_io_en),
    .io_out(r_count_6_io_out)
  );
  MyCounter r_count_7 ( // @[SWChisel.scala 171:41]
    .clock(r_count_7_clock),
    .reset(r_count_7_reset),
    .io_en(r_count_7_io_en),
    .io_out(r_count_7_io_out)
  );
  MyCounter r_count_8 ( // @[SWChisel.scala 171:41]
    .clock(r_count_8_clock),
    .reset(r_count_8_reset),
    .io_en(r_count_8_io_en),
    .io_out(r_count_8_io_out)
  );
  MyCounter r_count_9 ( // @[SWChisel.scala 171:41]
    .clock(r_count_9_clock),
    .reset(r_count_9_reset),
    .io_en(r_count_9_io_en),
    .io_out(r_count_9_io_out)
  );
  MAX max ( // @[SWChisel.scala 174:19]
    .clock(max_clock),
    .reset(max_reset),
    .io_start(max_io_start),
    .io_in(max_io_in),
    .io_done(max_io_done),
    .io_out(max_io_out)
  );
  assign io_result = max_io_out; // @[SWChisel.scala 181:13]
  assign io_done = max_io_done; // @[SWChisel.scala 182:11]
  assign array_0_io_q = io_q_0_b; // @[SWChisel.scala 220:19]
  assign array_0_io_r = 7'h63 == r_count_0_io_out ? io_r_99_b : _GEN_128; // @[SWChisel.scala 221:{19,19}]
  assign array_0_io_e_i = E_0; // @[SWChisel.scala 196:21]
  assign array_0_io_f_i = 16'sh0; // @[SWChisel.scala 198:21]
  assign array_0_io_ve_i = V1_1; // @[SWChisel.scala 197:22]
  assign array_0_io_vf_i = V1_0; // @[SWChisel.scala 199:22]
  assign array_0_io_vv_i = V2_0; // @[SWChisel.scala 200:22]
  assign array_1_io_q = io_q_1_b; // @[SWChisel.scala 220:19]
  assign array_1_io_r = 7'h63 == r_count_1_io_out ? io_r_99_b : _GEN_228; // @[SWChisel.scala 221:{19,19}]
  assign array_1_io_e_i = E_1; // @[SWChisel.scala 196:21]
  assign array_1_io_f_i = F_1; // @[SWChisel.scala 198:21]
  assign array_1_io_ve_i = V1_2; // @[SWChisel.scala 197:22]
  assign array_1_io_vf_i = V1_1; // @[SWChisel.scala 199:22]
  assign array_1_io_vv_i = V2_1; // @[SWChisel.scala 200:22]
  assign array_2_io_q = io_q_2_b; // @[SWChisel.scala 220:19]
  assign array_2_io_r = 7'h63 == r_count_2_io_out ? io_r_99_b : _GEN_328; // @[SWChisel.scala 221:{19,19}]
  assign array_2_io_e_i = E_2; // @[SWChisel.scala 196:21]
  assign array_2_io_f_i = F_2; // @[SWChisel.scala 198:21]
  assign array_2_io_ve_i = V1_3; // @[SWChisel.scala 197:22]
  assign array_2_io_vf_i = V1_2; // @[SWChisel.scala 199:22]
  assign array_2_io_vv_i = V2_2; // @[SWChisel.scala 200:22]
  assign array_3_io_q = io_q_3_b; // @[SWChisel.scala 220:19]
  assign array_3_io_r = 7'h63 == r_count_3_io_out ? io_r_99_b : _GEN_428; // @[SWChisel.scala 221:{19,19}]
  assign array_3_io_e_i = E_3; // @[SWChisel.scala 196:21]
  assign array_3_io_f_i = F_3; // @[SWChisel.scala 198:21]
  assign array_3_io_ve_i = V1_4; // @[SWChisel.scala 197:22]
  assign array_3_io_vf_i = V1_3; // @[SWChisel.scala 199:22]
  assign array_3_io_vv_i = V2_3; // @[SWChisel.scala 200:22]
  assign array_4_io_q = io_q_4_b; // @[SWChisel.scala 220:19]
  assign array_4_io_r = 7'h63 == r_count_4_io_out ? io_r_99_b : _GEN_528; // @[SWChisel.scala 221:{19,19}]
  assign array_4_io_e_i = E_4; // @[SWChisel.scala 196:21]
  assign array_4_io_f_i = F_4; // @[SWChisel.scala 198:21]
  assign array_4_io_ve_i = V1_5; // @[SWChisel.scala 197:22]
  assign array_4_io_vf_i = V1_4; // @[SWChisel.scala 199:22]
  assign array_4_io_vv_i = V2_4; // @[SWChisel.scala 200:22]
  assign array_5_io_q = io_q_5_b; // @[SWChisel.scala 220:19]
  assign array_5_io_r = 7'h63 == r_count_5_io_out ? io_r_99_b : _GEN_628; // @[SWChisel.scala 221:{19,19}]
  assign array_5_io_e_i = E_5; // @[SWChisel.scala 196:21]
  assign array_5_io_f_i = F_5; // @[SWChisel.scala 198:21]
  assign array_5_io_ve_i = V1_6; // @[SWChisel.scala 197:22]
  assign array_5_io_vf_i = V1_5; // @[SWChisel.scala 199:22]
  assign array_5_io_vv_i = V2_5; // @[SWChisel.scala 200:22]
  assign array_6_io_q = io_q_6_b; // @[SWChisel.scala 220:19]
  assign array_6_io_r = 7'h63 == r_count_6_io_out ? io_r_99_b : _GEN_728; // @[SWChisel.scala 221:{19,19}]
  assign array_6_io_e_i = E_6; // @[SWChisel.scala 196:21]
  assign array_6_io_f_i = F_6; // @[SWChisel.scala 198:21]
  assign array_6_io_ve_i = V1_7; // @[SWChisel.scala 197:22]
  assign array_6_io_vf_i = V1_6; // @[SWChisel.scala 199:22]
  assign array_6_io_vv_i = V2_6; // @[SWChisel.scala 200:22]
  assign array_7_io_q = io_q_7_b; // @[SWChisel.scala 220:19]
  assign array_7_io_r = 7'h63 == r_count_7_io_out ? io_r_99_b : _GEN_828; // @[SWChisel.scala 221:{19,19}]
  assign array_7_io_e_i = E_7; // @[SWChisel.scala 196:21]
  assign array_7_io_f_i = F_7; // @[SWChisel.scala 198:21]
  assign array_7_io_ve_i = V1_8; // @[SWChisel.scala 197:22]
  assign array_7_io_vf_i = V1_7; // @[SWChisel.scala 199:22]
  assign array_7_io_vv_i = V2_7; // @[SWChisel.scala 200:22]
  assign array_8_io_q = io_q_8_b; // @[SWChisel.scala 220:19]
  assign array_8_io_r = 7'h63 == r_count_8_io_out ? io_r_99_b : _GEN_928; // @[SWChisel.scala 221:{19,19}]
  assign array_8_io_e_i = E_8; // @[SWChisel.scala 196:21]
  assign array_8_io_f_i = F_8; // @[SWChisel.scala 198:21]
  assign array_8_io_ve_i = V1_9; // @[SWChisel.scala 197:22]
  assign array_8_io_vf_i = V1_8; // @[SWChisel.scala 199:22]
  assign array_8_io_vv_i = V2_8; // @[SWChisel.scala 200:22]
  assign array_9_io_q = io_q_9_b; // @[SWChisel.scala 220:19]
  assign array_9_io_r = 7'h63 == r_count_9_io_out ? io_r_99_b : _GEN_1028; // @[SWChisel.scala 221:{19,19}]
  assign array_9_io_e_i = E_9; // @[SWChisel.scala 196:21]
  assign array_9_io_f_i = F_9; // @[SWChisel.scala 198:21]
  assign array_9_io_ve_i = V1_10; // @[SWChisel.scala 197:22]
  assign array_9_io_vf_i = V1_9; // @[SWChisel.scala 199:22]
  assign array_9_io_vv_i = V2_9; // @[SWChisel.scala 200:22]
  assign r_count_0_clock = clock;
  assign r_count_0_reset = reset;
  assign r_count_0_io_en = start_reg_0; // @[SWChisel.scala 192:22]
  assign r_count_1_clock = clock;
  assign r_count_1_reset = reset;
  assign r_count_1_io_en = start_reg_1; // @[SWChisel.scala 192:22]
  assign r_count_2_clock = clock;
  assign r_count_2_reset = reset;
  assign r_count_2_io_en = start_reg_2; // @[SWChisel.scala 192:22]
  assign r_count_3_clock = clock;
  assign r_count_3_reset = reset;
  assign r_count_3_io_en = start_reg_3; // @[SWChisel.scala 192:22]
  assign r_count_4_clock = clock;
  assign r_count_4_reset = reset;
  assign r_count_4_io_en = start_reg_4; // @[SWChisel.scala 192:22]
  assign r_count_5_clock = clock;
  assign r_count_5_reset = reset;
  assign r_count_5_io_en = start_reg_5; // @[SWChisel.scala 192:22]
  assign r_count_6_clock = clock;
  assign r_count_6_reset = reset;
  assign r_count_6_io_en = start_reg_6; // @[SWChisel.scala 192:22]
  assign r_count_7_clock = clock;
  assign r_count_7_reset = reset;
  assign r_count_7_io_en = start_reg_7; // @[SWChisel.scala 192:22]
  assign r_count_8_clock = clock;
  assign r_count_8_reset = reset;
  assign r_count_8_io_en = start_reg_8; // @[SWChisel.scala 192:22]
  assign r_count_9_clock = clock;
  assign r_count_9_reset = reset;
  assign r_count_9_io_en = start_reg_9; // @[SWChisel.scala 192:22]
  assign max_clock = clock;
  assign max_reset = reset;
  assign max_io_start = start_reg_9; // @[SWChisel.scala 178:16]
  assign max_io_in = V1_10; // @[SWChisel.scala 177:13]
  always @(posedge clock) begin
    if (reset) begin // @[SWChisel.scala 162:18]
      E_0 <= -16'sh2; // @[SWChisel.scala 162:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      E_0 <= array_0_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_1 <= -16'sh3; // @[SWChisel.scala 162:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      E_1 <= array_1_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_2 <= -16'sh4; // @[SWChisel.scala 162:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      E_2 <= array_2_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_3 <= -16'sh5; // @[SWChisel.scala 162:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      E_3 <= array_3_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_4 <= -16'sh6; // @[SWChisel.scala 162:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      E_4 <= array_4_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_5 <= -16'sh7; // @[SWChisel.scala 162:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      E_5 <= array_5_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_6 <= -16'sh8; // @[SWChisel.scala 162:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      E_6 <= array_6_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_7 <= -16'sh9; // @[SWChisel.scala 162:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      E_7 <= array_7_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_8 <= -16'sha; // @[SWChisel.scala 162:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      E_8 <= array_8_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_9 <= -16'shb; // @[SWChisel.scala 162:18]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      E_9 <= array_9_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_1 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      F_1 <= array_0_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_2 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      F_2 <= array_1_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_3 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      F_3 <= array_2_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_4 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      F_4 <= array_3_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_5 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      F_5 <= array_4_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_6 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      F_6 <= array_5_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_7 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      F_7 <= array_6_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_8 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      F_8 <= array_7_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_9 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      F_9 <= array_8_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_0 <= -16'sh1; // @[SWChisel.scala 164:19]
    end else begin
      V1_0 <= 16'sh0; // @[SWChisel.scala 165:9]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_1 <= -16'sh2; // @[SWChisel.scala 164:19]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      V1_1 <= array_0_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_2 <= -16'sh3; // @[SWChisel.scala 164:19]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      V1_2 <= array_1_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_3 <= -16'sh4; // @[SWChisel.scala 164:19]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      V1_3 <= array_2_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_4 <= -16'sh5; // @[SWChisel.scala 164:19]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      V1_4 <= array_3_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_5 <= -16'sh6; // @[SWChisel.scala 164:19]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      V1_5 <= array_4_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_6 <= -16'sh7; // @[SWChisel.scala 164:19]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      V1_6 <= array_5_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_7 <= -16'sh8; // @[SWChisel.scala 164:19]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      V1_7 <= array_6_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_8 <= -16'sh9; // @[SWChisel.scala 164:19]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      V1_8 <= array_7_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_9 <= -16'sha; // @[SWChisel.scala 164:19]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      V1_9 <= array_8_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_10 <= -16'shb; // @[SWChisel.scala 164:19]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      V1_10 <= array_9_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_0 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_0 <= V1_0; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_1 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_1 <= V1_1; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_2 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_2 <= V1_2; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_3 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_3 <= V1_3; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_4 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_4 <= V1_4; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_5 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_5 <= V1_5; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_6 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_6 <= V1_6; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_7 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_7 <= V1_7; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_8 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_8 <= V1_8; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_9 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_9 <= V1_9; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_0 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_0 <= io_start; // @[SWChisel.scala 185:16]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_1 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_1 <= start_reg_0; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_2 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_2 <= start_reg_1; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_3 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_3 <= start_reg_2; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_4 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_4 <= start_reg_3; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_5 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_5 <= start_reg_4; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_6 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_6 <= start_reg_5; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_7 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_7 <= start_reg_6; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_8 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_8 <= start_reg_7; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_9 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_9 <= start_reg_8; // @[SWChisel.scala 187:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  E_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  E_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  E_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  E_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  E_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  E_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  E_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  E_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  E_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  E_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  F_1 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  F_2 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  F_3 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  F_4 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  F_5 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  F_6 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  F_7 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  F_8 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  F_9 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  V1_0 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  V1_1 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  V1_2 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  V1_3 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  V1_4 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  V1_5 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  V1_6 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  V1_7 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  V1_8 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  V1_9 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  V1_10 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  V2_0 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  V2_1 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  V2_2 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  V2_3 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  V2_4 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  V2_5 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  V2_6 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  V2_7 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  V2_8 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  V2_9 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  start_reg_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  start_reg_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  start_reg_2 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  start_reg_3 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  start_reg_4 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  start_reg_5 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  start_reg_6 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  start_reg_7 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  start_reg_8 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  start_reg_9 = _RAND_49[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
